// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.0.0 Build 614 04/24/2018 SJ Standard Edition"

// DATE "01/19/2026 15:17:20"

// 
// Device: Altera EP4CE15F17C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module fftsign (
	clk,
	reset_n,
	sink_valid,
	sink_ready,
	sink_error,
	sink_sop,
	sink_eop,
	sink_real,
	sink_imag,
	inverse,
	source_valid,
	source_ready,
	source_error,
	source_sop,
	source_eop,
	source_real,
	source_imag,
	source_exp)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	sink_valid;
output 	sink_ready;
input 	[1:0] sink_error;
input 	sink_sop;
input 	sink_eop;
input 	[9:0] sink_real;
input 	[9:0] sink_imag;
input 	[0:0] inverse;
output 	source_valid;
input 	source_ready;
output 	[1:0] source_error;
output 	source_sop;
output 	source_eop;
output 	[9:0] source_real;
output 	[9:0] source_imag;
output 	[5:0] source_exp;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;
wire \~GND~combout ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \source_ready~input_o ;
wire \sink_valid~input_o ;
wire \sink_eop~input_o ;
wire \sink_sop~input_o ;
wire \sink_error[0]~input_o ;
wire \sink_error[1]~input_o ;
wire \inverse[0]~input_o ;
wire \sink_imag[2]~input_o ;
wire \sink_real[2]~input_o ;
wire \sink_imag[1]~input_o ;
wire \sink_real[1]~input_o ;
wire \sink_imag[0]~input_o ;
wire \sink_real[0]~input_o ;
wire \sink_imag[9]~input_o ;
wire \sink_real[9]~input_o ;
wire \sink_imag[8]~input_o ;
wire \sink_real[8]~input_o ;
wire \sink_imag[7]~input_o ;
wire \sink_real[7]~input_o ;
wire \sink_imag[6]~input_o ;
wire \sink_real[6]~input_o ;
wire \sink_imag[5]~input_o ;
wire \sink_real[5]~input_o ;
wire \sink_imag[4]~input_o ;
wire \sink_real[4]~input_o ;
wire \sink_imag[3]~input_o ;
wire \sink_real[3]~input_o ;


fftsign_fftsign_fft_ii_0 fft_ii_0(
	.at_sink_ready_s(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ),
	.at_source_valid_s(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ),
	.at_source_error_0(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ),
	.at_source_error_1(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ),
	.at_source_sop_s(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ),
	.at_source_eop_s(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ),
	.at_source_data_16(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ),
	.at_source_data_17(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ),
	.at_source_data_18(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ),
	.at_source_data_19(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ),
	.at_source_data_20(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ),
	.at_source_data_21(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ),
	.at_source_data_22(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ),
	.at_source_data_23(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ),
	.at_source_data_24(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ),
	.at_source_data_25(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ),
	.at_source_data_6(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ),
	.at_source_data_7(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ),
	.at_source_data_8(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ),
	.at_source_data_9(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ),
	.at_source_data_10(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ),
	.at_source_data_11(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ),
	.at_source_data_12(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ),
	.at_source_data_13(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ),
	.at_source_data_14(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ),
	.at_source_data_15(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ),
	.at_source_data_0(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ),
	.at_source_data_1(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ),
	.at_source_data_2(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ),
	.at_source_data_3(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ),
	.at_source_data_4(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ),
	.at_source_data_5(\fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ),
	.GND_port(\~GND~combout ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.source_ready(\source_ready~input_o ),
	.sink_valid(\sink_valid~input_o ),
	.sink_eop(\sink_eop~input_o ),
	.sink_sop(\sink_sop~input_o ),
	.sink_error_0(\sink_error[0]~input_o ),
	.sink_error_1(\sink_error[1]~input_o ),
	.inverse_0(\inverse[0]~input_o ),
	.sink_imag_2(\sink_imag[2]~input_o ),
	.sink_real_2(\sink_real[2]~input_o ),
	.sink_imag_1(\sink_imag[1]~input_o ),
	.sink_real_1(\sink_real[1]~input_o ),
	.sink_imag_0(\sink_imag[0]~input_o ),
	.sink_real_0(\sink_real[0]~input_o ),
	.sink_imag_9(\sink_imag[9]~input_o ),
	.sink_real_9(\sink_real[9]~input_o ),
	.sink_imag_8(\sink_imag[8]~input_o ),
	.sink_real_8(\sink_real[8]~input_o ),
	.sink_imag_7(\sink_imag[7]~input_o ),
	.sink_real_7(\sink_real[7]~input_o ),
	.sink_imag_6(\sink_imag[6]~input_o ),
	.sink_real_6(\sink_real[6]~input_o ),
	.sink_imag_5(\sink_imag[5]~input_o ),
	.sink_real_5(\sink_real[5]~input_o ),
	.sink_imag_4(\sink_imag[4]~input_o ),
	.sink_real_4(\sink_real[4]~input_o ),
	.sink_imag_3(\sink_imag[3]~input_o ),
	.sink_real_3(\sink_real[3]~input_o ));

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \source_ready~input_o  = source_ready;

assign \sink_valid~input_o  = sink_valid;

assign \sink_eop~input_o  = sink_eop;

assign \sink_sop~input_o  = sink_sop;

assign \sink_error[0]~input_o  = sink_error[0];

assign \sink_error[1]~input_o  = sink_error[1];

assign \inverse[0]~input_o  = inverse[0];

assign \sink_imag[2]~input_o  = sink_imag[2];

assign \sink_real[2]~input_o  = sink_real[2];

assign \sink_imag[1]~input_o  = sink_imag[1];

assign \sink_real[1]~input_o  = sink_real[1];

assign \sink_imag[0]~input_o  = sink_imag[0];

assign \sink_real[0]~input_o  = sink_real[0];

assign \sink_imag[9]~input_o  = sink_imag[9];

assign \sink_real[9]~input_o  = sink_real[9];

assign \sink_imag[8]~input_o  = sink_imag[8];

assign \sink_real[8]~input_o  = sink_real[8];

assign \sink_imag[7]~input_o  = sink_imag[7];

assign \sink_real[7]~input_o  = sink_real[7];

assign \sink_imag[6]~input_o  = sink_imag[6];

assign \sink_real[6]~input_o  = sink_real[6];

assign \sink_imag[5]~input_o  = sink_imag[5];

assign \sink_real[5]~input_o  = sink_real[5];

assign \sink_imag[4]~input_o  = sink_imag[4];

assign \sink_real[4]~input_o  = sink_real[4];

assign \sink_imag[3]~input_o  = sink_imag[3];

assign \sink_real[3]~input_o  = sink_real[3];

assign sink_ready = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;

assign source_valid = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;

assign source_error[0] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;

assign source_error[1] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;

assign source_sop = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;

assign source_eop = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;

assign source_real[0] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;

assign source_real[1] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;

assign source_real[2] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;

assign source_real[3] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;

assign source_real[4] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;

assign source_real[5] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;

assign source_real[6] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[22]~q ;

assign source_real[7] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[23]~q ;

assign source_real[8] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[24]~q ;

assign source_real[9] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[25]~q ;

assign source_imag[0] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;

assign source_imag[1] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;

assign source_imag[2] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;

assign source_imag[3] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;

assign source_imag[4] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;

assign source_imag[5] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;

assign source_imag[6] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;

assign source_imag[7] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;

assign source_imag[8] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;

assign source_imag[9] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;

assign source_exp[0] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;

assign source_exp[1] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;

assign source_exp[2] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;

assign source_exp[3] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;

assign source_exp[4] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;

assign source_exp[5] = \fft_ii_0|asj_fft_si_se_so_b_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;

endmodule

module fftsign_fftsign_fft_ii_0 (
	at_sink_ready_s,
	at_source_valid_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_22,
	at_source_data_23,
	at_source_data_24,
	at_source_data_25,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_14,
	at_source_data_15,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	GND_port,
	clk,
	reset_n,
	source_ready,
	sink_valid,
	sink_eop,
	sink_sop,
	sink_error_0,
	sink_error_1,
	inverse_0,
	sink_imag_2,
	sink_real_2,
	sink_imag_1,
	sink_real_1,
	sink_imag_0,
	sink_real_0,
	sink_imag_9,
	sink_real_9,
	sink_imag_8,
	sink_real_8,
	sink_imag_7,
	sink_real_7,
	sink_imag_6,
	sink_real_6,
	sink_imag_5,
	sink_real_5,
	sink_imag_4,
	sink_real_4,
	sink_imag_3,
	sink_real_3)/* synthesis synthesis_greybox=1 */;
output 	at_sink_ready_s;
output 	at_source_valid_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_22;
output 	at_source_data_23;
output 	at_source_data_24;
output 	at_source_data_25;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_valid;
input 	sink_eop;
input 	sink_sop;
input 	sink_error_0;
input 	sink_error_1;
input 	inverse_0;
input 	sink_imag_2;
input 	sink_real_2;
input 	sink_imag_1;
input 	sink_real_1;
input 	sink_imag_0;
input 	sink_real_0;
input 	sink_imag_9;
input 	sink_real_9;
input 	sink_imag_8;
input 	sink_real_8;
input 	sink_imag_7;
input 	sink_real_7;
input 	sink_imag_6;
input 	sink_real_6;
input 	sink_imag_5;
input 	sink_real_5;
input 	sink_imag_4;
input 	sink_real_4;
input 	sink_imag_3;
input 	sink_real_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_asj_fft_si_se_so_b asj_fft_si_se_so_b_inst(
	.at_sink_ready_s(at_sink_ready_s),
	.at_source_valid_s(at_source_valid_s),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s(at_source_sop_s),
	.at_source_eop_s(at_source_eop_s),
	.at_source_data_16(at_source_data_16),
	.at_source_data_17(at_source_data_17),
	.at_source_data_18(at_source_data_18),
	.at_source_data_19(at_source_data_19),
	.at_source_data_20(at_source_data_20),
	.at_source_data_21(at_source_data_21),
	.at_source_data_22(at_source_data_22),
	.at_source_data_23(at_source_data_23),
	.at_source_data_24(at_source_data_24),
	.at_source_data_25(at_source_data_25),
	.at_source_data_6(at_source_data_6),
	.at_source_data_7(at_source_data_7),
	.at_source_data_8(at_source_data_8),
	.at_source_data_9(at_source_data_9),
	.at_source_data_10(at_source_data_10),
	.at_source_data_11(at_source_data_11),
	.at_source_data_12(at_source_data_12),
	.at_source_data_13(at_source_data_13),
	.at_source_data_14(at_source_data_14),
	.at_source_data_15(at_source_data_15),
	.at_source_data_0(at_source_data_0),
	.at_source_data_1(at_source_data_1),
	.at_source_data_2(at_source_data_2),
	.at_source_data_3(at_source_data_3),
	.at_source_data_4(at_source_data_4),
	.at_source_data_5(at_source_data_5),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready),
	.sink_valid(sink_valid),
	.sink_eop(sink_eop),
	.sink_sop(sink_sop),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.inverse_0(inverse_0),
	.sink_imag({sink_imag_9,sink_imag_8,sink_imag_7,sink_imag_6,sink_imag_5,sink_imag_4,sink_imag_3,sink_imag_2,sink_imag_1,sink_imag_0}),
	.sink_real({sink_real_9,sink_real_8,sink_real_7,sink_real_6,sink_real_5,sink_real_4,sink_real_3,sink_real_2,sink_real_1,sink_real_0}));

endmodule

module fftsign_asj_fft_si_se_so_b (
	at_sink_ready_s,
	at_source_valid_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_22,
	at_source_data_23,
	at_source_data_24,
	at_source_data_25,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_14,
	at_source_data_15,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	GND_port,
	clk,
	reset_n,
	source_ready,
	sink_valid,
	sink_eop,
	sink_sop,
	sink_error_0,
	sink_error_1,
	inverse_0,
	sink_imag,
	sink_real)/* synthesis synthesis_greybox=1 */;
output 	at_sink_ready_s;
output 	at_source_valid_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_22;
output 	at_source_data_23;
output 	at_source_data_24;
output 	at_source_data_25;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_valid;
input 	sink_eop;
input 	sink_sop;
input 	sink_error_0;
input 	sink_error_1;
input 	inverse_0;
input 	[9:0] sink_imag;
input 	[9:0] sink_real;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \master_sink_ena~q ;
wire \sink_in_work~q ;
wire \data_count_sig[7]~q ;
wire \data_count_sig[9]~q ;
wire \data_count_sig[8]~q ;
wire \data_count_sig[3]~q ;
wire \data_count_sig[4]~q ;
wire \data_count_sig[6]~q ;
wire \data_count_sig[5]~q ;
wire \data_count_sig[2]~q ;
wire \data_count_sig[0]~q ;
wire \data_count_sig[1]~q ;
wire \data_count_sig[0]~11 ;
wire \data_count_sig[0]~10_combout ;
wire \data_count_sig[1]~13 ;
wire \data_count_sig[1]~12_combout ;
wire \data_count_sig[2]~15 ;
wire \data_count_sig[2]~14_combout ;
wire \data_count_sig[3]~17 ;
wire \data_count_sig[3]~16_combout ;
wire \data_count_sig[4]~19 ;
wire \data_count_sig[4]~18_combout ;
wire \data_count_sig[5]~21 ;
wire \data_count_sig[5]~20_combout ;
wire \data_count_sig[6]~23 ;
wire \data_count_sig[6]~22_combout ;
wire \data_count_sig[7]~25 ;
wire \data_count_sig[7]~24_combout ;
wire \data_count_sig[8]~30 ;
wire \data_count_sig[8]~29_combout ;
wire \data_count_sig[9]~31_combout ;
wire \writer|rdy_for_next_block~q ;
wire \writer|disable_wr~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][9]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][8]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \sel_we|lpp_c_i~q ;
wire \writer|data_rdy_int~q ;
wire \writer|wren[3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][2]~q ;
wire \ram_cxb_wr|ram_in_reg[3][1]~q ;
wire \ram_cxb_wr|ram_in_reg[3][3]~q ;
wire \ram_cxb_wr|ram_in_reg[3][5]~q ;
wire \ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ;
wire \ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ;
wire \writer|wren[0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][2]~q ;
wire \ram_cxb_wr|ram_in_reg[0][1]~q ;
wire \ram_cxb_wr|ram_in_reg[0][3]~q ;
wire \ram_cxb_wr|ram_in_reg[0][5]~q ;
wire \writer|wren[1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][2]~q ;
wire \ram_cxb_wr|ram_in_reg[1][1]~q ;
wire \ram_cxb_wr|ram_in_reg[1][3]~q ;
wire \ram_cxb_wr|ram_in_reg[1][5]~q ;
wire \writer|wren[2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][2]~q ;
wire \ram_cxb_wr|ram_in_reg[2][1]~q ;
wire \ram_cxb_wr|ram_in_reg[2][3]~q ;
wire \ram_cxb_wr|ram_in_reg[2][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][9]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][8]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][3]~q ;
wire \ctrl|blk_done_int~q ;
wire \get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ;
wire \get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ;
wire \core_real_in[2]~q ;
wire \core_imag_in[2]~q ;
wire \core_real_in[1]~q ;
wire \core_imag_in[1]~q ;
wire \core_real_in[0]~q ;
wire \core_imag_in[0]~q ;
wire \core_real_in[9]~q ;
wire \core_imag_in[9]~q ;
wire \core_real_in[8]~q ;
wire \core_imag_in[8]~q ;
wire \core_real_in[7]~q ;
wire \core_imag_in[7]~q ;
wire \core_real_in[6]~q ;
wire \core_imag_in[6]~q ;
wire \core_real_in[5]~q ;
wire \core_imag_in[5]~q ;
wire \core_real_in[4]~q ;
wire \core_imag_in[4]~q ;
wire \core_real_in[3]~q ;
wire \core_imag_in[3]~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2~portbdataout ;
wire \twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3~portbdataout ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ;
wire \twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ;
wire \twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ;
wire \ram_cxb_bfp_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][8]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][9]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][9]~q ;
wire \auk_dsp_interface_controller_1|source_packet_error[1]~q ;
wire \auk_dsp_interface_controller_1|source_packet_error[0]~q ;
wire \auk_dsp_interface_controller_1|source_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_stall_reg~q ;
wire \auk_dsp_atlantic_sink_1|send_eop_s~q ;
wire \auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ;
wire \auk_dsp_atlantic_sink_1|sink_start~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ;
wire \auk_dsp_atlantic_sink_1|sink_stall~combout ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[1]~q ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[0]~q ;
wire \master_source_ena~q ;
wire \sink_ready_ctrl_d~q ;
wire \auk_dsp_atlantic_sink_1|send_sop_s~q ;
wire \sop~q ;
wire \global_clock_enable~0_combout ;
wire \auk_dsp_interface_controller_1|stall_reg~q ;
wire \auk_dsp_atlantic_source_1|source_stall_int_d~q ;
wire \fft_real_out[0]~q ;
wire \fft_real_out[1]~q ;
wire \fft_real_out[2]~q ;
wire \fft_real_out[3]~q ;
wire \fft_real_out[4]~q ;
wire \fft_real_out[5]~q ;
wire \fft_real_out[6]~q ;
wire \fft_real_out[7]~q ;
wire \fft_real_out[8]~q ;
wire \fft_real_out[9]~q ;
wire \fft_imag_out[0]~q ;
wire \fft_imag_out[1]~q ;
wire \fft_imag_out[2]~q ;
wire \fft_imag_out[3]~q ;
wire \fft_imag_out[4]~q ;
wire \fft_imag_out[5]~q ;
wire \fft_imag_out[6]~q ;
wire \fft_imag_out[7]~q ;
wire \fft_imag_out[8]~q ;
wire \fft_imag_out[9]~q ;
wire \exponent_out[0]~q ;
wire \exponent_out[1]~q ;
wire \exponent_out[2]~q ;
wire \exponent_out[3]~q ;
wire \exponent_out[4]~q ;
wire \exponent_out[5]~q ;
wire \auk_dsp_atlantic_source_1|Mux0~1_combout ;
wire \fft_s1_cur.WAIT_FOR_INPUT~q ;
wire \fft_s1_cur.WRITE_INPUT~q ;
wire \fft_s1_cur.IDLE~q ;
wire \WideOr1~0_combout ;
wire \global_clock_enable~1_combout ;
wire \sink_in_work~0_combout ;
wire \val_out~q ;
wire \oe~q ;
wire \master_source_ena~0_combout ;
wire \sop~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \master_source_sop~q ;
wire \data_count_sig[9]~26_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \data_count_sig[9]~27_combout ;
wire \data_count_sig[3]~28_combout ;
wire \exponent_out[2]~0_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[0]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[0]~q ;
wire \fft_dirn~q ;
wire \fft_real_out~0_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[1]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[1]~q ;
wire \fft_real_out~1_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[2]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[2]~q ;
wire \fft_real_out~2_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[3]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[3]~q ;
wire \fft_real_out~3_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[4]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[4]~q ;
wire \fft_real_out~4_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[5]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[5]~q ;
wire \fft_real_out~5_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[6]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[6]~q ;
wire \fft_real_out~6_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[7]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[7]~q ;
wire \fft_real_out~7_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[8]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[8]~q ;
wire \fft_real_out~8_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[9]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[9]~q ;
wire \fft_real_out~9_combout ;
wire \fft_imag_out~0_combout ;
wire \fft_imag_out~1_combout ;
wire \fft_imag_out~2_combout ;
wire \fft_imag_out~3_combout ;
wire \fft_imag_out~4_combout ;
wire \fft_imag_out~5_combout ;
wire \fft_imag_out~6_combout ;
wire \fft_imag_out~7_combout ;
wire \fft_imag_out~8_combout ;
wire \fft_imag_out~9_combout ;
wire \bfpc|blk_exp[0]~q ;
wire \exponent_out~1_combout ;
wire \bfpc|blk_exp[1]~q ;
wire \exponent_out~2_combout ;
wire \bfpc|blk_exp[2]~q ;
wire \exponent_out~3_combout ;
wire \bfpc|blk_exp[3]~q ;
wire \exponent_out~4_combout ;
wire \bfpc|blk_exp[4]~q ;
wire \exponent_out~5_combout ;
wire \bfpc|blk_exp[5]~q ;
wire \exponent_out~6_combout ;
wire \fft_s1_cur.NO_WRITE~q ;
wire \fft_s1_cur.DONE_WRITING~q ;
wire \fft_s1_cur.EARLY_DONE~q ;
wire \fft_s1_cur.WAIT_FOR_INPUT~0_combout ;
wire \fft_s1_cur.FFT_PROCESS_A~q ;
wire \fft_s1_cur.WAIT_FOR_INPUT~1_combout ;
wire \eop_out~q ;
wire \data_rdy_vec[24]~q ;
wire \fft_s1_cur.NO_WRITE~0_combout ;
wire \no_del_input_blk:delay_next_block|tdl_arr[0]~q ;
wire \fft_s1_cur.NO_WRITE~1_combout ;
wire \fft_s1_cur.NO_WRITE~2_combout ;
wire \fft_s1_cur.NO_WRITE~3_combout ;
wire \fft_s1_cur.WAIT_FOR_INPUT~2_combout ;
wire \fft_s1_cur.WRITE_INPUT~0_combout ;
wire \fft_s1_cur.NO_WRITE~4_combout ;
wire \fft_s1_cur.WAIT_FOR_INPUT~3_combout ;
wire \fft_s2_cur.START_LPP~q ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~q ;
wire \bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ;
wire \val_out~0_combout ;
wire \fft_s2_cur.LPP_OUTPUT_RDY~q ;
wire \fft_s2_cur.LPP_DONE~q ;
wire \val_out~1_combout ;
wire \sop_out~q ;
wire \master_source_sop~0_combout ;
wire \sel_we|wait_count[0]~0_combout ;
wire \inv_i~q ;
wire \fft_dirn~0_combout ;
wire \exp_en~q ;
wire \fft_s1_cur.NO_WRITE~5_combout ;
wire \fft_s1_cur.DONE_WRITING~0_combout ;
wire \fft_s1_cur.EARLY_DONE~0_combout ;
wire \fft_s1_cur.FFT_PROCESS_A~0_combout ;
wire \eop_out~0_combout ;
wire \data_rdy_vec[23]~q ;
wire \data_rdy_vec~0_combout ;
wire \gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ;
wire \fft_s2_cur.START_LPP~0_combout ;
wire \gen_radix_4_last_pass:lpp|gen_burst_val:delay_val|tdl_arr[4]~q ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~0_combout ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~1_combout ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~2_combout ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~3_combout ;
wire \fft_s2_cur.LPP_OUTPUT_RDY~0_combout ;
wire \fft_s2_cur.LPP_DONE~0_combout ;
wire \delay_sop|tdl_arr[6]~q ;
wire \sop_out~0_combout ;
wire \sop_out~1_combout ;
wire \sop_out~2_combout ;
wire \inv_i~0_combout ;
wire \bfpc|slb_last[0]~q ;
wire \bfpc|slb_last[1]~q ;
wire \bfpc|slb_last[2]~q ;
wire \data_rdy_vec[22]~q ;
wire \data_rdy_vec~1_combout ;
wire \bfpdft|gen_disc:bfp_detect|slb_i[0]~q ;
wire \bfpdft|gen_disc:bfp_detect|slb_i[1]~q ;
wire \bfpdft|gen_disc:bfp_detect|slb_i[2]~q ;
wire \bfpdft|gen_disc:bfp_detect|slb_i[3]~q ;
wire \bfpdft|gen_disc:bfp_detect|Mux2~0_combout ;
wire \delay_blk_done|tdl_arr[23]~q ;
wire \bfpdft|gen_disc:bfp_detect|Mux1~0_combout ;
wire \data_rdy_vec[21]~q ;
wire \data_rdy_vec~2_combout ;
wire \bfpc|gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[6]~q ;
wire \data_rdy_vec[20]~q ;
wire \data_rdy_vec~3_combout ;
wire \bfpdft|reg_no_twiddle[6][0][5]~q ;
wire \bfpdft|reg_no_twiddle[6][0][9]~q ;
wire \bfpdft|reg_no_twiddle[6][1][5]~q ;
wire \bfpdft|reg_no_twiddle[6][1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ;
wire \bfpdft|reg_no_twiddle[6][0][6]~q ;
wire \bfpdft|reg_no_twiddle[6][1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ;
wire \bfpdft|reg_no_twiddle[6][0][7]~q ;
wire \bfpdft|reg_no_twiddle[6][1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ;
wire \bfpdft|reg_no_twiddle[6][0][8]~q ;
wire \bfpdft|reg_no_twiddle[6][1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ;
wire \data_rdy_vec[19]~q ;
wire \data_rdy_vec~4_combout ;
wire \lpp_ram_data_out[3][12]~q ;
wire \lpp_ram_data_out[0][12]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ;
wire \lpp_ram_data_out[1][12]~q ;
wire \lpp_ram_data_out[2][12]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ;
wire \lpp_ram_data_out[3][2]~q ;
wire \lpp_ram_data_out[0][2]~q ;
wire \lpp_ram_data_out[1][2]~q ;
wire \lpp_ram_data_out[2][2]~q ;
wire \lpp_ram_data_out[3][11]~q ;
wire \lpp_ram_data_out[0][11]~q ;
wire \lpp_ram_data_out[1][11]~q ;
wire \lpp_ram_data_out[2][11]~q ;
wire \lpp_ram_data_out[3][1]~q ;
wire \lpp_ram_data_out[0][1]~q ;
wire \lpp_ram_data_out[1][1]~q ;
wire \lpp_ram_data_out[2][1]~q ;
wire \lpp_ram_data_out[3][10]~q ;
wire \lpp_ram_data_out[0][10]~q ;
wire \lpp_ram_data_out[1][10]~q ;
wire \lpp_ram_data_out[2][10]~q ;
wire \lpp_ram_data_out[3][0]~q ;
wire \lpp_ram_data_out[0][0]~q ;
wire \lpp_ram_data_out[1][0]~q ;
wire \lpp_ram_data_out[2][0]~q ;
wire \lpp_ram_data_out[3][19]~q ;
wire \lpp_ram_data_out[0][19]~q ;
wire \lpp_ram_data_out[1][19]~q ;
wire \lpp_ram_data_out[2][19]~q ;
wire \lpp_ram_data_out[3][9]~q ;
wire \lpp_ram_data_out[0][9]~q ;
wire \lpp_ram_data_out[1][9]~q ;
wire \lpp_ram_data_out[2][9]~q ;
wire \lpp_ram_data_out[3][18]~q ;
wire \lpp_ram_data_out[0][18]~q ;
wire \lpp_ram_data_out[1][18]~q ;
wire \lpp_ram_data_out[2][18]~q ;
wire \lpp_ram_data_out[3][8]~q ;
wire \lpp_ram_data_out[0][8]~q ;
wire \lpp_ram_data_out[1][8]~q ;
wire \lpp_ram_data_out[2][8]~q ;
wire \lpp_ram_data_out[3][17]~q ;
wire \lpp_ram_data_out[0][17]~q ;
wire \lpp_ram_data_out[1][17]~q ;
wire \lpp_ram_data_out[2][17]~q ;
wire \lpp_ram_data_out[3][7]~q ;
wire \lpp_ram_data_out[0][7]~q ;
wire \lpp_ram_data_out[1][7]~q ;
wire \lpp_ram_data_out[2][7]~q ;
wire \lpp_ram_data_out[3][16]~q ;
wire \lpp_ram_data_out[0][16]~q ;
wire \lpp_ram_data_out[1][16]~q ;
wire \lpp_ram_data_out[2][16]~q ;
wire \lpp_ram_data_out[3][6]~q ;
wire \lpp_ram_data_out[0][6]~q ;
wire \lpp_ram_data_out[1][6]~q ;
wire \lpp_ram_data_out[2][6]~q ;
wire \lpp_ram_data_out[3][15]~q ;
wire \lpp_ram_data_out[0][15]~q ;
wire \lpp_ram_data_out[1][15]~q ;
wire \lpp_ram_data_out[2][15]~q ;
wire \lpp_ram_data_out[3][5]~q ;
wire \lpp_ram_data_out[0][5]~q ;
wire \lpp_ram_data_out[1][5]~q ;
wire \lpp_ram_data_out[2][5]~q ;
wire \lpp_ram_data_out[3][14]~q ;
wire \lpp_ram_data_out[0][14]~q ;
wire \lpp_ram_data_out[1][14]~q ;
wire \lpp_ram_data_out[2][14]~q ;
wire \lpp_ram_data_out[3][4]~q ;
wire \lpp_ram_data_out[0][4]~q ;
wire \lpp_ram_data_out[1][4]~q ;
wire \lpp_ram_data_out[2][4]~q ;
wire \lpp_ram_data_out[3][13]~q ;
wire \lpp_ram_data_out[0][13]~q ;
wire \lpp_ram_data_out[1][13]~q ;
wire \lpp_ram_data_out[2][13]~q ;
wire \lpp_ram_data_out[3][3]~q ;
wire \lpp_ram_data_out[0][3]~q ;
wire \lpp_ram_data_out[1][3]~q ;
wire \lpp_ram_data_out[2][3]~q ;
wire \data_rdy_vec[18]~q ;
wire \data_rdy_vec~5_combout ;
wire \lpp_c_en_vec[6]~q ;
wire \lpp_c_en_vec[1]~q ;
wire \lpp_ram_data_out~0_combout ;
wire \lpp_ram_data_out~1_combout ;
wire \lpp_ram_data_out~2_combout ;
wire \lpp_ram_data_out~3_combout ;
wire \lpp_ram_data_out~4_combout ;
wire \lpp_ram_data_out~5_combout ;
wire \lpp_ram_data_out~6_combout ;
wire \lpp_ram_data_out~7_combout ;
wire \lpp_ram_data_out~8_combout ;
wire \lpp_ram_data_out~9_combout ;
wire \lpp_ram_data_out~10_combout ;
wire \lpp_ram_data_out~11_combout ;
wire \lpp_ram_data_out~12_combout ;
wire \lpp_ram_data_out~13_combout ;
wire \lpp_ram_data_out~14_combout ;
wire \lpp_ram_data_out~15_combout ;
wire \lpp_ram_data_out~16_combout ;
wire \lpp_ram_data_out~17_combout ;
wire \lpp_ram_data_out~18_combout ;
wire \lpp_ram_data_out~19_combout ;
wire \lpp_ram_data_out~20_combout ;
wire \lpp_ram_data_out~21_combout ;
wire \lpp_ram_data_out~22_combout ;
wire \lpp_ram_data_out~23_combout ;
wire \lpp_ram_data_out~24_combout ;
wire \lpp_ram_data_out~25_combout ;
wire \lpp_ram_data_out~26_combout ;
wire \lpp_ram_data_out~27_combout ;
wire \lpp_ram_data_out~28_combout ;
wire \lpp_ram_data_out~29_combout ;
wire \lpp_ram_data_out~30_combout ;
wire \lpp_ram_data_out~31_combout ;
wire \lpp_ram_data_out~32_combout ;
wire \lpp_ram_data_out~33_combout ;
wire \lpp_ram_data_out~34_combout ;
wire \lpp_ram_data_out~35_combout ;
wire \lpp_ram_data_out~36_combout ;
wire \lpp_ram_data_out~37_combout ;
wire \lpp_ram_data_out~38_combout ;
wire \lpp_ram_data_out~39_combout ;
wire \lpp_ram_data_out~40_combout ;
wire \lpp_ram_data_out~41_combout ;
wire \lpp_ram_data_out~42_combout ;
wire \lpp_ram_data_out~43_combout ;
wire \lpp_ram_data_out~44_combout ;
wire \lpp_ram_data_out~45_combout ;
wire \lpp_ram_data_out~46_combout ;
wire \lpp_ram_data_out~47_combout ;
wire \lpp_ram_data_out~48_combout ;
wire \lpp_ram_data_out~49_combout ;
wire \lpp_ram_data_out~50_combout ;
wire \lpp_ram_data_out~51_combout ;
wire \lpp_ram_data_out~52_combout ;
wire \lpp_ram_data_out~53_combout ;
wire \lpp_ram_data_out~54_combout ;
wire \lpp_ram_data_out~55_combout ;
wire \lpp_ram_data_out~56_combout ;
wire \lpp_ram_data_out~57_combout ;
wire \lpp_ram_data_out~58_combout ;
wire \lpp_ram_data_out~59_combout ;
wire \lpp_ram_data_out~60_combout ;
wire \lpp_ram_data_out~61_combout ;
wire \lpp_ram_data_out~62_combout ;
wire \lpp_ram_data_out~63_combout ;
wire \lpp_ram_data_out~64_combout ;
wire \lpp_ram_data_out~65_combout ;
wire \lpp_ram_data_out~66_combout ;
wire \lpp_ram_data_out~67_combout ;
wire \lpp_ram_data_out~68_combout ;
wire \lpp_ram_data_out~69_combout ;
wire \lpp_ram_data_out~70_combout ;
wire \lpp_ram_data_out~71_combout ;
wire \lpp_ram_data_out~72_combout ;
wire \lpp_ram_data_out~73_combout ;
wire \lpp_ram_data_out~74_combout ;
wire \lpp_ram_data_out~75_combout ;
wire \lpp_ram_data_out~76_combout ;
wire \lpp_ram_data_out~77_combout ;
wire \lpp_ram_data_out~78_combout ;
wire \lpp_ram_data_out~79_combout ;
wire \data_rdy_vec[17]~q ;
wire \data_rdy_vec~6_combout ;
wire \gen_radix_4_last_pass:gen_lpp_addr|en_d~q ;
wire \wren_a[3]~q ;
wire \ccc|a_ram_data_in_bus[12]~q ;
wire \ccc|wraddress_a_bus[0]~q ;
wire \ccc|wraddress_a_bus[1]~q ;
wire \ccc|wraddress_a_bus[18]~q ;
wire \ccc|wraddress_a_bus[3]~q ;
wire \ccc|wraddress_a_bus[20]~q ;
wire \ccc|wraddress_a_bus[5]~q ;
wire \ccc|wraddress_a_bus[14]~q ;
wire \ccc|wraddress_a_bus[15]~q ;
wire \ccc|rdaddress_a_bus[0]~q ;
wire \ccc|rdaddress_a_bus[1]~q ;
wire \ccc|rdaddress_a_bus[18]~q ;
wire \ccc|rdaddress_a_bus[3]~q ;
wire \ccc|rdaddress_a_bus[20]~q ;
wire \ccc|rdaddress_a_bus[5]~q ;
wire \ccc|rdaddress_a_bus[22]~q ;
wire \ccc|rdaddress_a_bus[7]~q ;
wire \lpp_c_en_vec[5]~q ;
wire \lpp_c_en_vec~0_combout ;
wire \lpp_c_en_vec~1_combout ;
wire \wren_a[0]~q ;
wire \ccc|a_ram_data_in_bus[72]~q ;
wire \ccc|wraddress_a_bus[24]~q ;
wire \ccc|wraddress_a_bus[25]~q ;
wire \ccc|wraddress_a_bus[10]~q ;
wire \ccc|wraddress_a_bus[27]~q ;
wire \ccc|wraddress_a_bus[12]~q ;
wire \ccc|wraddress_a_bus[29]~q ;
wire \ccc|rdaddress_a_bus[24]~q ;
wire \ccc|rdaddress_a_bus[25]~q ;
wire \ccc|rdaddress_a_bus[10]~q ;
wire \ccc|rdaddress_a_bus[27]~q ;
wire \ccc|rdaddress_a_bus[12]~q ;
wire \ccc|rdaddress_a_bus[29]~q ;
wire \ccc|rdaddress_a_bus[14]~q ;
wire \ccc|rdaddress_a_bus[31]~q ;
wire \wren_a[1]~q ;
wire \ccc|a_ram_data_in_bus[52]~q ;
wire \ccc|wraddress_a_bus[17]~q ;
wire \ccc|wraddress_a_bus[19]~q ;
wire \ccc|wraddress_a_bus[21]~q ;
wire \ccc|rdaddress_a_bus[17]~q ;
wire \ccc|rdaddress_a_bus[19]~q ;
wire \ccc|rdaddress_a_bus[21]~q ;
wire \ccc|rdaddress_a_bus[23]~q ;
wire \wren_a[2]~q ;
wire \ccc|a_ram_data_in_bus[32]~q ;
wire \ccc|wraddress_a_bus[9]~q ;
wire \ccc|wraddress_a_bus[11]~q ;
wire \ccc|wraddress_a_bus[13]~q ;
wire \ccc|rdaddress_a_bus[9]~q ;
wire \ccc|rdaddress_a_bus[11]~q ;
wire \ccc|rdaddress_a_bus[13]~q ;
wire \ccc|rdaddress_a_bus[15]~q ;
wire \ccc|a_ram_data_in_bus[2]~q ;
wire \ccc|a_ram_data_in_bus[62]~q ;
wire \ccc|a_ram_data_in_bus[42]~q ;
wire \ccc|a_ram_data_in_bus[22]~q ;
wire \ccc|a_ram_data_in_bus[11]~q ;
wire \ccc|a_ram_data_in_bus[71]~q ;
wire \ccc|a_ram_data_in_bus[51]~q ;
wire \ccc|a_ram_data_in_bus[31]~q ;
wire \ccc|a_ram_data_in_bus[1]~q ;
wire \ccc|a_ram_data_in_bus[61]~q ;
wire \ccc|a_ram_data_in_bus[41]~q ;
wire \ccc|a_ram_data_in_bus[21]~q ;
wire \ccc|a_ram_data_in_bus[10]~q ;
wire \ccc|a_ram_data_in_bus[70]~q ;
wire \ccc|a_ram_data_in_bus[50]~q ;
wire \ccc|a_ram_data_in_bus[30]~q ;
wire \ccc|a_ram_data_in_bus[0]~q ;
wire \ccc|a_ram_data_in_bus[60]~q ;
wire \ccc|a_ram_data_in_bus[40]~q ;
wire \ccc|a_ram_data_in_bus[20]~q ;
wire \ccc|a_ram_data_in_bus[19]~q ;
wire \ccc|a_ram_data_in_bus[79]~q ;
wire \ccc|a_ram_data_in_bus[59]~q ;
wire \ccc|a_ram_data_in_bus[39]~q ;
wire \ccc|a_ram_data_in_bus[9]~q ;
wire \ccc|a_ram_data_in_bus[69]~q ;
wire \ccc|a_ram_data_in_bus[49]~q ;
wire \ccc|a_ram_data_in_bus[29]~q ;
wire \ccc|a_ram_data_in_bus[18]~q ;
wire \ccc|a_ram_data_in_bus[78]~q ;
wire \ccc|a_ram_data_in_bus[58]~q ;
wire \ccc|a_ram_data_in_bus[38]~q ;
wire \ccc|a_ram_data_in_bus[8]~q ;
wire \ccc|a_ram_data_in_bus[68]~q ;
wire \ccc|a_ram_data_in_bus[48]~q ;
wire \ccc|a_ram_data_in_bus[28]~q ;
wire \ccc|a_ram_data_in_bus[17]~q ;
wire \ccc|a_ram_data_in_bus[77]~q ;
wire \ccc|a_ram_data_in_bus[57]~q ;
wire \ccc|a_ram_data_in_bus[37]~q ;
wire \ccc|a_ram_data_in_bus[7]~q ;
wire \ccc|a_ram_data_in_bus[67]~q ;
wire \ccc|a_ram_data_in_bus[47]~q ;
wire \ccc|a_ram_data_in_bus[27]~q ;
wire \ccc|a_ram_data_in_bus[16]~q ;
wire \ccc|a_ram_data_in_bus[76]~q ;
wire \ccc|a_ram_data_in_bus[56]~q ;
wire \ccc|a_ram_data_in_bus[36]~q ;
wire \ccc|a_ram_data_in_bus[6]~q ;
wire \ccc|a_ram_data_in_bus[66]~q ;
wire \ccc|a_ram_data_in_bus[46]~q ;
wire \ccc|a_ram_data_in_bus[26]~q ;
wire \ccc|a_ram_data_in_bus[15]~q ;
wire \ccc|a_ram_data_in_bus[75]~q ;
wire \ccc|a_ram_data_in_bus[55]~q ;
wire \ccc|a_ram_data_in_bus[35]~q ;
wire \ccc|a_ram_data_in_bus[5]~q ;
wire \ccc|a_ram_data_in_bus[65]~q ;
wire \ccc|a_ram_data_in_bus[45]~q ;
wire \ccc|a_ram_data_in_bus[25]~q ;
wire \ccc|a_ram_data_in_bus[14]~q ;
wire \ccc|a_ram_data_in_bus[74]~q ;
wire \ccc|a_ram_data_in_bus[54]~q ;
wire \ccc|a_ram_data_in_bus[34]~q ;
wire \ccc|a_ram_data_in_bus[4]~q ;
wire \ccc|a_ram_data_in_bus[64]~q ;
wire \ccc|a_ram_data_in_bus[44]~q ;
wire \ccc|a_ram_data_in_bus[24]~q ;
wire \ccc|a_ram_data_in_bus[13]~q ;
wire \ccc|a_ram_data_in_bus[73]~q ;
wire \ccc|a_ram_data_in_bus[53]~q ;
wire \ccc|a_ram_data_in_bus[33]~q ;
wire \ccc|a_ram_data_in_bus[3]~q ;
wire \ccc|a_ram_data_in_bus[63]~q ;
wire \ccc|a_ram_data_in_bus[43]~q ;
wire \ccc|a_ram_data_in_bus[23]~q ;
wire \data_rdy_vec[16]~q ;
wire \data_rdy_vec~7_combout ;
wire \sel_we|wc_i_d~q ;
wire \wc_vec[3]~q ;
wire \wren_a~2_combout ;
wire \fft_s1_cur.WAIT_FOR_INPUT~4_combout ;
wire \wren_a~3_combout ;
wire \writer|data_in_r[2]~q ;
wire \sel_ram_in~q ;
wire \ram_cxb_wr|ram_in_reg[1][0]~q ;
wire \writer|wr_address_i_int[0]~q ;
wire \data_rdy_vec[2]~q ;
wire \writer|wr_address_i_int[1]~q ;
wire \ram_cxb_wr|ram_in_reg[1][2]~q ;
wire \writer|wr_address_i_int[2]~q ;
wire \writer|wr_address_i_int[3]~q ;
wire \ram_cxb_wr|ram_in_reg[1][4]~q ;
wire \writer|wr_address_i_int[4]~q ;
wire \writer|wr_address_i_int[5]~q ;
wire \writer|wr_address_i_int[6]~q ;
wire \writer|wr_address_i_int[7]~q ;
wire \ram_cxb_rd|ram_in_reg[1][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ;
wire \data_rdy_vec[0]~q ;
wire \ram_cxb_rd|ram_in_reg[3][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ;
wire \ram_cxb_rd|ram_in_reg[1][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ;
wire \ram_cxb_rd|ram_in_reg[3][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ;
wire \ram_cxb_rd|ram_in_reg[1][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ;
wire \ram_cxb_rd|ram_in_reg[3][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ;
wire \ram_cxb_rd|ram_in_reg[0][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ;
wire \ram_cxb_rd|ram_in_reg[0][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[3][7]~q ;
wire \lpp_c_en_vec[4]~q ;
wire \lpp_c_en_vec~2_combout ;
wire \wren_a~4_combout ;
wire \ram_cxb_wr|ram_in_reg[0][0]~q ;
wire \ram_cxb_wr|ram_in_reg[0][2]~q ;
wire \ram_cxb_wr|ram_in_reg[0][4]~q ;
wire \ram_cxb_rd|ram_in_reg[0][0]~q ;
wire \ram_cxb_rd|ram_in_reg[0][1]~q ;
wire \ram_cxb_rd|ram_in_reg[0][2]~q ;
wire \ram_cxb_rd|ram_in_reg[0][3]~q ;
wire \ram_cxb_rd|ram_in_reg[0][4]~q ;
wire \ram_cxb_rd|ram_in_reg[0][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[2][7]~q ;
wire \wren_a~5_combout ;
wire \ram_cxb_rd|ram_in_reg[1][1]~q ;
wire \ram_cxb_rd|ram_in_reg[1][3]~q ;
wire \ram_cxb_rd|ram_in_reg[1][5]~q ;
wire \wren_a~6_combout ;
wire \ram_cxb_rd|ram_in_reg[2][1]~q ;
wire \ram_cxb_rd|ram_in_reg[2][3]~q ;
wire \ram_cxb_rd|ram_in_reg[2][5]~q ;
wire \writer|data_in_i[2]~q ;
wire \writer|data_in_r[1]~q ;
wire \writer|data_in_i[1]~q ;
wire \writer|data_in_r[0]~q ;
wire \writer|data_in_i[0]~q ;
wire \writer|data_in_r[9]~q ;
wire \writer|data_in_i[9]~q ;
wire \writer|data_in_r[8]~q ;
wire \writer|data_in_i[8]~q ;
wire \writer|data_in_r[7]~q ;
wire \writer|data_in_i[7]~q ;
wire \writer|data_in_r[6]~q ;
wire \writer|data_in_i[6]~q ;
wire \writer|data_in_r[5]~q ;
wire \writer|data_in_i[5]~q ;
wire \writer|data_in_r[4]~q ;
wire \writer|data_in_i[4]~q ;
wire \writer|data_in_r[3]~q ;
wire \writer|data_in_i[3]~q ;
wire \data_rdy_vec[15]~q ;
wire \data_rdy_vec~8_combout ;
wire \wc_vec[2]~q ;
wire \wc_vec~0_combout ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ;
wire \bfpdft|reg_no_twiddle[6][0][2]~q ;
wire \sel_ram_in~0_combout ;
wire \get_wr_swtiches|swa_tdl[16][0]~q ;
wire \data_rdy_vec[1]~q ;
wire \data_rdy_vec~9_combout ;
wire \get_wr_swtiches|swa_tdl[16][1]~q ;
wire \rd_adgen|rd_addr_c[0]~q ;
wire \rd_adgen|rd_addr_d[0]~q ;
wire \rd_adgen|sw[0]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ;
wire \data_rdy_vec~10_combout ;
wire \rd_adgen|rd_addr_b[1]~q ;
wire \rd_adgen|rd_addr_d[1]~q ;
wire \rd_adgen|sw[1]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ;
wire \rd_adgen|rd_addr_c[2]~q ;
wire \rd_adgen|rd_addr_d[2]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[2]~q ;
wire \rd_adgen|rd_addr_b[3]~q ;
wire \rd_adgen|rd_addr_d[3]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[3]~q ;
wire \rd_adgen|rd_addr_c[4]~q ;
wire \rd_adgen|rd_addr_d[4]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[4]~q ;
wire \rd_adgen|rd_addr_b[5]~q ;
wire \rd_adgen|rd_addr_d[5]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[5]~q ;
wire \rd_adgen|rd_addr_d[6]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ;
wire \rd_adgen|rd_addr_d[7]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ;
wire \lpp_c_en_vec[3]~q ;
wire \lpp_c_en_vec~3_combout ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ;
wire \bfpdft|reg_no_twiddle[6][1][2]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ;
wire \bfpdft|reg_no_twiddle[6][0][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ;
wire \bfpdft|reg_no_twiddle[6][1][1]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ;
wire \bfpdft|reg_no_twiddle[6][0][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ;
wire \bfpdft|reg_no_twiddle[6][1][0]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ;
wire \bfpdft|reg_no_twiddle[6][0][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ;
wire \bfpdft|reg_no_twiddle[6][1][4]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ;
wire \bfpdft|reg_no_twiddle[6][0][3]~q ;
wire \bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ;
wire \bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ;
wire \bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ;
wire \bfpdft|reg_no_twiddle[6][1][3]~q ;
wire \data_rdy_vec[14]~q ;
wire \data_rdy_vec~11_combout ;
wire \p_cd_en[2]~q ;
wire \wc_vec[1]~q ;
wire \wc_vec~1_combout ;
wire \ctrl|p[2]~q ;
wire \ctrl|p[0]~q ;
wire \ctrl|p[1]~q ;
wire \ctrl|k_count[4]~q ;
wire \ctrl|k_count[0]~q ;
wire \ctrl|k_count[2]~q ;
wire \rd_adgen|Add1~0_combout ;
wire \rd_adgen|Mux1~0_combout ;
wire \rd_adgen|Mux1~1_combout ;
wire \ctrl|k_count[6]~q ;
wire \ctrl|k_count[1]~q ;
wire \ctrl|k_count[3]~q ;
wire \rd_adgen|Add0~0_combout ;
wire \ctrl|k_count[5]~q ;
wire \rd_adgen|Add1~1_combout ;
wire \rd_adgen|Add1~2_combout ;
wire \rd_adgen|Mux0~0_combout ;
wire \rd_adgen|Mux0~1_combout ;
wire \ctrl|k_count[7]~q ;
wire \data_imag_in_reg[2]~q ;
wire \data_real_in_reg[2]~q ;
wire \core_real_in~0_combout ;
wire \data_rdy_vec~12_combout ;
wire \twid_factors|Mux0~0_combout ;
wire \lpp_c_en_vec[2]~q ;
wire \lpp_c_en_vec~4_combout ;
wire \core_imag_in~0_combout ;
wire \data_imag_in_reg[1]~q ;
wire \data_real_in_reg[1]~q ;
wire \core_real_in~1_combout ;
wire \core_imag_in~1_combout ;
wire \data_imag_in_reg[0]~q ;
wire \data_real_in_reg[0]~q ;
wire \core_real_in~2_combout ;
wire \core_imag_in~2_combout ;
wire \data_imag_in_reg[9]~q ;
wire \data_real_in_reg[9]~q ;
wire \core_real_in~3_combout ;
wire \core_imag_in~3_combout ;
wire \data_imag_in_reg[8]~q ;
wire \data_real_in_reg[8]~q ;
wire \core_real_in~4_combout ;
wire \core_imag_in~4_combout ;
wire \data_imag_in_reg[7]~q ;
wire \data_real_in_reg[7]~q ;
wire \core_real_in~5_combout ;
wire \core_imag_in~5_combout ;
wire \data_imag_in_reg[6]~q ;
wire \data_real_in_reg[6]~q ;
wire \core_real_in~6_combout ;
wire \core_imag_in~6_combout ;
wire \data_imag_in_reg[5]~q ;
wire \data_real_in_reg[5]~q ;
wire \core_real_in~7_combout ;
wire \core_imag_in~7_combout ;
wire \data_imag_in_reg[4]~q ;
wire \data_real_in_reg[4]~q ;
wire \core_real_in~8_combout ;
wire \core_imag_in~8_combout ;
wire \data_imag_in_reg[3]~q ;
wire \data_real_in_reg[3]~q ;
wire \core_real_in~9_combout ;
wire \core_imag_in~9_combout ;
wire \delay_np|tdl_arr[9]~q ;
wire \data_rdy_vec[13]~q ;
wire \data_rdy_vec~13_combout ;
wire \p_tdl[13][2]~q ;
wire \p_tdl[13][0]~q ;
wire \p_tdl[13][1]~q ;
wire \p_tdl[11][0]~q ;
wire \reg_we_window~0_combout ;
wire \p_tdl[11][2]~q ;
wire \p_tdl[11][1]~q ;
wire \reg_we_window~1_combout ;
wire \wc_vec~2_combout ;
wire \data_rdy_vec[4]~q ;
wire \ctrl|next_pass_i~q ;
wire \data_imag_in_reg~0_combout ;
wire \data_real_in_reg~0_combout ;
wire \lpp_c_en_vec~5_combout ;
wire \data_imag_in_reg~1_combout ;
wire \data_real_in_reg~1_combout ;
wire \data_imag_in_reg~2_combout ;
wire \data_real_in_reg~2_combout ;
wire \data_imag_in_reg~3_combout ;
wire \data_real_in_reg~3_combout ;
wire \data_imag_in_reg~4_combout ;
wire \data_real_in_reg~4_combout ;
wire \data_imag_in_reg~5_combout ;
wire \data_real_in_reg~5_combout ;
wire \data_imag_in_reg~6_combout ;
wire \data_real_in_reg~6_combout ;
wire \data_imag_in_reg~7_combout ;
wire \data_real_in_reg~7_combout ;
wire \data_imag_in_reg~8_combout ;
wire \data_real_in_reg~8_combout ;
wire \data_imag_in_reg~9_combout ;
wire \data_real_in_reg~9_combout ;
wire \twiddle_data[0][1][0]~q ;
wire \twiddle_data[0][1][1]~q ;
wire \twiddle_data[0][1][2]~q ;
wire \twiddle_data[0][1][3]~q ;
wire \twiddle_data[0][1][4]~q ;
wire \twiddle_data[0][1][5]~q ;
wire \twiddle_data[0][1][6]~q ;
wire \twiddle_data[0][1][7]~q ;
wire \twiddle_data[0][1][8]~q ;
wire \twiddle_data[0][1][9]~q ;
wire \twiddle_data[0][0][0]~q ;
wire \twiddle_data[0][0][1]~q ;
wire \twiddle_data[0][0][2]~q ;
wire \twiddle_data[0][0][3]~q ;
wire \twiddle_data[0][0][4]~q ;
wire \twiddle_data[0][0][5]~q ;
wire \twiddle_data[0][0][6]~q ;
wire \twiddle_data[0][0][7]~q ;
wire \twiddle_data[0][0][8]~q ;
wire \twiddle_data[0][0][9]~q ;
wire \twiddle_data[1][1][0]~q ;
wire \twiddle_data[1][1][1]~q ;
wire \twiddle_data[1][1][2]~q ;
wire \twiddle_data[1][1][3]~q ;
wire \twiddle_data[1][1][4]~q ;
wire \twiddle_data[1][1][5]~q ;
wire \twiddle_data[1][1][6]~q ;
wire \twiddle_data[1][1][7]~q ;
wire \twiddle_data[1][1][8]~q ;
wire \twiddle_data[1][1][9]~q ;
wire \twiddle_data[1][0][0]~q ;
wire \twiddle_data[1][0][1]~q ;
wire \twiddle_data[1][0][2]~q ;
wire \twiddle_data[1][0][3]~q ;
wire \twiddle_data[1][0][4]~q ;
wire \twiddle_data[1][0][5]~q ;
wire \twiddle_data[1][0][6]~q ;
wire \twiddle_data[1][0][7]~q ;
wire \twiddle_data[1][0][8]~q ;
wire \twiddle_data[1][0][9]~q ;
wire \twiddle_data[2][1][0]~q ;
wire \twiddle_data[2][1][1]~q ;
wire \twiddle_data[2][1][2]~q ;
wire \twiddle_data[2][1][3]~q ;
wire \twiddle_data[2][1][4]~q ;
wire \twiddle_data[2][1][5]~q ;
wire \twiddle_data[2][1][6]~q ;
wire \twiddle_data[2][1][7]~q ;
wire \twiddle_data[2][1][8]~q ;
wire \twiddle_data[2][1][9]~q ;
wire \twiddle_data[2][0][0]~q ;
wire \twiddle_data[2][0][1]~q ;
wire \twiddle_data[2][0][2]~q ;
wire \twiddle_data[2][0][3]~q ;
wire \twiddle_data[2][0][4]~q ;
wire \twiddle_data[2][0][5]~q ;
wire \twiddle_data[2][0][6]~q ;
wire \twiddle_data[2][0][7]~q ;
wire \twiddle_data[2][0][8]~q ;
wire \twiddle_data[2][0][9]~q ;
wire \data_rdy_vec[12]~q ;
wire \data_rdy_vec~14_combout ;
wire \p_tdl[12][2]~q ;
wire \p_tdl~0_combout ;
wire \p_tdl[12][0]~q ;
wire \p_tdl~1_combout ;
wire \p_tdl[12][1]~q ;
wire \p_tdl~2_combout ;
wire \p_tdl[10][0]~q ;
wire \p_tdl~3_combout ;
wire \p_tdl[10][2]~q ;
wire \p_tdl~4_combout ;
wire \p_tdl[10][1]~q ;
wire \p_tdl~5_combout ;
wire \data_rdy_vec[3]~q ;
wire \data_rdy_vec~15_combout ;
wire \twiddle_data~0_combout ;
wire \twiddle_data~1_combout ;
wire \twiddle_data~2_combout ;
wire \twiddle_data~3_combout ;
wire \twiddle_data~4_combout ;
wire \twiddle_data~5_combout ;
wire \twiddle_data~6_combout ;
wire \twiddle_data~7_combout ;
wire \twiddle_data~8_combout ;
wire \twiddle_data~9_combout ;
wire \twiddle_data~10_combout ;
wire \twiddle_data~11_combout ;
wire \twiddle_data~12_combout ;
wire \twiddle_data~13_combout ;
wire \twiddle_data~14_combout ;
wire \twiddle_data~15_combout ;
wire \twiddle_data~16_combout ;
wire \twiddle_data~17_combout ;
wire \twiddle_data~18_combout ;
wire \twiddle_data~19_combout ;
wire \twiddle_data~20_combout ;
wire \twiddle_data~21_combout ;
wire \twiddle_data~22_combout ;
wire \twiddle_data~23_combout ;
wire \twiddle_data~24_combout ;
wire \twiddle_data~25_combout ;
wire \twiddle_data~26_combout ;
wire \twiddle_data~27_combout ;
wire \twiddle_data~28_combout ;
wire \twiddle_data~29_combout ;
wire \twiddle_data~30_combout ;
wire \twiddle_data~31_combout ;
wire \twiddle_data~32_combout ;
wire \twiddle_data~33_combout ;
wire \twiddle_data~34_combout ;
wire \twiddle_data~35_combout ;
wire \twiddle_data~36_combout ;
wire \twiddle_data~37_combout ;
wire \twiddle_data~38_combout ;
wire \twiddle_data~39_combout ;
wire \twiddle_data~40_combout ;
wire \twiddle_data~41_combout ;
wire \twiddle_data~42_combout ;
wire \twiddle_data~43_combout ;
wire \twiddle_data~44_combout ;
wire \twiddle_data~45_combout ;
wire \twiddle_data~46_combout ;
wire \twiddle_data~47_combout ;
wire \twiddle_data~48_combout ;
wire \twiddle_data~49_combout ;
wire \twiddle_data~50_combout ;
wire \twiddle_data~51_combout ;
wire \twiddle_data~52_combout ;
wire \twiddle_data~53_combout ;
wire \twiddle_data~54_combout ;
wire \twiddle_data~55_combout ;
wire \twiddle_data~56_combout ;
wire \twiddle_data~57_combout ;
wire \twiddle_data~58_combout ;
wire \twiddle_data~59_combout ;
wire \data_rdy_vec[11]~q ;
wire \data_rdy_vec~16_combout ;
wire \p_tdl~6_combout ;
wire \p_tdl~7_combout ;
wire \p_tdl~8_combout ;
wire \p_tdl[9][0]~q ;
wire \p_tdl~9_combout ;
wire \p_tdl[9][2]~q ;
wire \p_tdl~10_combout ;
wire \p_tdl[9][1]~q ;
wire \p_tdl~11_combout ;
wire \data_rdy_vec~17_combout ;
wire \rd_adgen|Mux1~5_combout ;
wire \rd_adgen|Mux1~6_combout ;
wire \rd_adgen|Mux0~5_combout ;
wire \rd_adgen|Mux0~6_combout ;
wire \data_rdy_vec[10]~q ;
wire \data_rdy_vec~18_combout ;
wire \p_tdl[8][0]~q ;
wire \p_tdl~12_combout ;
wire \p_tdl[8][2]~q ;
wire \p_tdl~13_combout ;
wire \p_tdl[8][1]~q ;
wire \p_tdl~14_combout ;
wire \data_rdy_vec[9]~q ;
wire \data_rdy_vec~19_combout ;
wire \p_tdl[7][0]~q ;
wire \p_tdl~15_combout ;
wire \p_tdl[7][2]~q ;
wire \p_tdl~16_combout ;
wire \p_tdl[7][1]~q ;
wire \p_tdl~17_combout ;
wire \data_rdy_vec[8]~q ;
wire \data_rdy_vec~20_combout ;
wire \p_tdl[6][0]~q ;
wire \p_tdl~18_combout ;
wire \p_tdl[6][2]~q ;
wire \p_tdl~19_combout ;
wire \p_tdl[6][1]~q ;
wire \p_tdl~20_combout ;
wire \ccc|ram_data_out0[17]~q ;
wire \ccc|ram_data_out1[17]~q ;
wire \sw_r_tdl[4][0]~q ;
wire \ccc|ram_data_out2[17]~q ;
wire \ccc|ram_data_out3[17]~q ;
wire \sw_r_tdl[4][1]~q ;
wire \ccc|ram_data_out0[15]~q ;
wire \ccc|ram_data_out1[15]~q ;
wire \ccc|ram_data_out2[15]~q ;
wire \ccc|ram_data_out3[15]~q ;
wire \ccc|ram_data_out0[16]~q ;
wire \ccc|ram_data_out1[16]~q ;
wire \ccc|ram_data_out2[16]~q ;
wire \ccc|ram_data_out3[16]~q ;
wire \ccc|ram_data_out0[18]~q ;
wire \ccc|ram_data_out1[18]~q ;
wire \ccc|ram_data_out2[18]~q ;
wire \ccc|ram_data_out3[18]~q ;
wire \ccc|ram_data_out0[14]~q ;
wire \ccc|ram_data_out1[14]~q ;
wire \ccc|ram_data_out2[14]~q ;
wire \ccc|ram_data_out3[14]~q ;
wire \ccc|ram_data_out2[13]~q ;
wire \ccc|ram_data_out3[13]~q ;
wire \ccc|ram_data_out0[13]~q ;
wire \ccc|ram_data_out1[13]~q ;
wire \ccc|ram_data_out2[12]~q ;
wire \ccc|ram_data_out3[12]~q ;
wire \ccc|ram_data_out0[12]~q ;
wire \ccc|ram_data_out1[12]~q ;
wire \ccc|ram_data_out2[11]~q ;
wire \ccc|ram_data_out3[11]~q ;
wire \ccc|ram_data_out0[11]~q ;
wire \ccc|ram_data_out1[11]~q ;
wire \ccc|ram_data_out2[10]~q ;
wire \ccc|ram_data_out3[10]~q ;
wire \ccc|ram_data_out0[10]~q ;
wire \ccc|ram_data_out1[10]~q ;
wire \ccc|ram_data_out0[19]~q ;
wire \ccc|ram_data_out1[19]~q ;
wire \ccc|ram_data_out2[19]~q ;
wire \ccc|ram_data_out3[19]~q ;
wire \ccc|ram_data_out0[5]~q ;
wire \ccc|ram_data_out1[5]~q ;
wire \ccc|ram_data_out2[5]~q ;
wire \ccc|ram_data_out3[5]~q ;
wire \ccc|ram_data_out0[6]~q ;
wire \ccc|ram_data_out1[6]~q ;
wire \ccc|ram_data_out2[6]~q ;
wire \ccc|ram_data_out3[6]~q ;
wire \ccc|ram_data_out0[7]~q ;
wire \ccc|ram_data_out1[7]~q ;
wire \ccc|ram_data_out2[7]~q ;
wire \ccc|ram_data_out3[7]~q ;
wire \ccc|ram_data_out0[8]~q ;
wire \ccc|ram_data_out1[8]~q ;
wire \ccc|ram_data_out2[8]~q ;
wire \ccc|ram_data_out3[8]~q ;
wire \ccc|ram_data_out0[4]~q ;
wire \ccc|ram_data_out1[4]~q ;
wire \ccc|ram_data_out2[4]~q ;
wire \ccc|ram_data_out3[4]~q ;
wire \ccc|ram_data_out2[3]~q ;
wire \ccc|ram_data_out3[3]~q ;
wire \ccc|ram_data_out0[3]~q ;
wire \ccc|ram_data_out1[3]~q ;
wire \ccc|ram_data_out2[2]~q ;
wire \ccc|ram_data_out3[2]~q ;
wire \ccc|ram_data_out0[2]~q ;
wire \ccc|ram_data_out1[2]~q ;
wire \ccc|ram_data_out2[1]~q ;
wire \ccc|ram_data_out3[1]~q ;
wire \ccc|ram_data_out0[1]~q ;
wire \ccc|ram_data_out1[1]~q ;
wire \ccc|ram_data_out2[0]~q ;
wire \ccc|ram_data_out3[0]~q ;
wire \ccc|ram_data_out0[0]~q ;
wire \ccc|ram_data_out1[0]~q ;
wire \ccc|ram_data_out0[9]~q ;
wire \ccc|ram_data_out1[9]~q ;
wire \ccc|ram_data_out2[9]~q ;
wire \ccc|ram_data_out3[9]~q ;
wire \data_rdy_vec[7]~q ;
wire \data_rdy_vec~21_combout ;
wire \p_tdl[5][0]~q ;
wire \p_tdl~21_combout ;
wire \p_tdl[5][2]~q ;
wire \p_tdl~22_combout ;
wire \p_tdl[5][1]~q ;
wire \p_tdl~23_combout ;
wire \sw_r_tdl[3][0]~q ;
wire \sw_r_tdl[3][1]~q ;
wire \data_rdy_vec[6]~q ;
wire \data_rdy_vec~22_combout ;
wire \p_tdl[4][0]~q ;
wire \p_tdl~24_combout ;
wire \p_tdl[4][2]~q ;
wire \p_tdl~25_combout ;
wire \p_tdl[4][1]~q ;
wire \p_tdl~26_combout ;
wire \sw_r_tdl[2][0]~q ;
wire \sw_r_tdl[2][1]~q ;
wire \data_rdy_vec[5]~q ;
wire \data_rdy_vec~23_combout ;
wire \p_tdl[3][0]~q ;
wire \p_tdl~27_combout ;
wire \p_tdl[3][2]~q ;
wire \p_tdl~28_combout ;
wire \p_tdl[3][1]~q ;
wire \p_tdl~29_combout ;
wire \sw_r_tdl[1][0]~q ;
wire \sw_r_tdl[1][1]~q ;
wire \data_rdy_vec~24_combout ;
wire \p_tdl[2][0]~q ;
wire \p_tdl~30_combout ;
wire \p_tdl[2][2]~q ;
wire \p_tdl~31_combout ;
wire \p_tdl[2][1]~q ;
wire \p_tdl~32_combout ;
wire \sw_r_tdl[0][0]~q ;
wire \sw_r_tdl[0][1]~q ;
wire \p_tdl[1][0]~q ;
wire \p_tdl~33_combout ;
wire \p_tdl[1][2]~q ;
wire \p_tdl~34_combout ;
wire \p_tdl[1][1]~q ;
wire \p_tdl~35_combout ;
wire \p_tdl[0][0]~q ;
wire \p_tdl~36_combout ;
wire \p_tdl[0][2]~q ;
wire \p_tdl~37_combout ;
wire \p_tdl[0][1]~q ;
wire \p_tdl~38_combout ;
wire \p_tdl~39_combout ;
wire \p_tdl~40_combout ;
wire \p_tdl~41_combout ;


fftsign_asj_fft_dft_bfp bfpdft(
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_8_0(\ram_cxb_bfp_data|ram_in_reg[0][8]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_8_2(\ram_cxb_bfp_data|ram_in_reg[2][8]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_8_1(\ram_cxb_bfp_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_8_3(\ram_cxb_bfp_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_9_0(\ram_cxb_bfp_data|ram_in_reg[0][9]~q ),
	.ram_in_reg_9_2(\ram_cxb_bfp_data|ram_in_reg[2][9]~q ),
	.ram_in_reg_9_1(\ram_cxb_bfp_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_3(\ram_cxb_bfp_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_8_4(\ram_cxb_bfp_data|ram_in_reg[4][8]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_8_6(\ram_cxb_bfp_data|ram_in_reg[6][8]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_8_5(\ram_cxb_bfp_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_8_7(\ram_cxb_bfp_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_9_4(\ram_cxb_bfp_data|ram_in_reg[4][9]~q ),
	.ram_in_reg_9_6(\ram_cxb_bfp_data|ram_in_reg[6][9]~q ),
	.ram_in_reg_9_5(\ram_cxb_bfp_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_9_7(\ram_cxb_bfp_data|ram_in_reg[7][9]~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_0(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.sdetdIDLE(\bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ),
	.slb_last_0(\bfpc|slb_last[0]~q ),
	.slb_last_1(\bfpc|slb_last[1]~q ),
	.slb_last_2(\bfpc|slb_last[2]~q ),
	.slb_i_0(\bfpdft|gen_disc:bfp_detect|slb_i[0]~q ),
	.slb_i_1(\bfpdft|gen_disc:bfp_detect|slb_i[1]~q ),
	.slb_i_2(\bfpdft|gen_disc:bfp_detect|slb_i[2]~q ),
	.slb_i_3(\bfpdft|gen_disc:bfp_detect|slb_i[3]~q ),
	.Mux2(\bfpdft|gen_disc:bfp_detect|Mux2~0_combout ),
	.Mux1(\bfpdft|gen_disc:bfp_detect|Mux1~0_combout ),
	.tdl_arr_6(\bfpc|gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[6]~q ),
	.reg_no_twiddle605(\bfpdft|reg_no_twiddle[6][0][5]~q ),
	.reg_no_twiddle609(\bfpdft|reg_no_twiddle[6][0][9]~q ),
	.reg_no_twiddle615(\bfpdft|reg_no_twiddle[6][1][5]~q ),
	.reg_no_twiddle619(\bfpdft|reg_no_twiddle[6][1][9]~q ),
	.tdl_arr_5_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.reg_no_twiddle606(\bfpdft|reg_no_twiddle[6][0][6]~q ),
	.reg_no_twiddle616(\bfpdft|reg_no_twiddle[6][1][6]~q ),
	.tdl_arr_6_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.reg_no_twiddle607(\bfpdft|reg_no_twiddle[6][0][7]~q ),
	.reg_no_twiddle617(\bfpdft|reg_no_twiddle[6][1][7]~q ),
	.tdl_arr_7_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.reg_no_twiddle608(\bfpdft|reg_no_twiddle[6][0][8]~q ),
	.reg_no_twiddle618(\bfpdft|reg_no_twiddle[6][1][8]~q ),
	.tdl_arr_8_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_2_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.reg_no_twiddle602(\bfpdft|reg_no_twiddle[6][0][2]~q ),
	.tdl_arr_2_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.reg_no_twiddle612(\bfpdft|reg_no_twiddle[6][1][2]~q ),
	.tdl_arr_1_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.reg_no_twiddle601(\bfpdft|reg_no_twiddle[6][0][1]~q ),
	.tdl_arr_1_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.reg_no_twiddle611(\bfpdft|reg_no_twiddle[6][1][1]~q ),
	.tdl_arr_0_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.reg_no_twiddle600(\bfpdft|reg_no_twiddle[6][0][0]~q ),
	.tdl_arr_0_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.reg_no_twiddle610(\bfpdft|reg_no_twiddle[6][1][0]~q ),
	.tdl_arr_4_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.reg_no_twiddle604(\bfpdft|reg_no_twiddle[6][0][4]~q ),
	.tdl_arr_4_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.reg_no_twiddle614(\bfpdft|reg_no_twiddle[6][1][4]~q ),
	.tdl_arr_3_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.reg_no_twiddle603(\bfpdft|reg_no_twiddle[6][0][3]~q ),
	.tdl_arr_3_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.reg_no_twiddle613(\bfpdft|reg_no_twiddle[6][1][3]~q ),
	.twiddle_data010(\twiddle_data[0][1][0]~q ),
	.twiddle_data011(\twiddle_data[0][1][1]~q ),
	.twiddle_data012(\twiddle_data[0][1][2]~q ),
	.twiddle_data013(\twiddle_data[0][1][3]~q ),
	.twiddle_data014(\twiddle_data[0][1][4]~q ),
	.twiddle_data015(\twiddle_data[0][1][5]~q ),
	.twiddle_data016(\twiddle_data[0][1][6]~q ),
	.twiddle_data017(\twiddle_data[0][1][7]~q ),
	.twiddle_data018(\twiddle_data[0][1][8]~q ),
	.twiddle_data019(\twiddle_data[0][1][9]~q ),
	.twiddle_data000(\twiddle_data[0][0][0]~q ),
	.twiddle_data001(\twiddle_data[0][0][1]~q ),
	.twiddle_data002(\twiddle_data[0][0][2]~q ),
	.twiddle_data003(\twiddle_data[0][0][3]~q ),
	.twiddle_data004(\twiddle_data[0][0][4]~q ),
	.twiddle_data005(\twiddle_data[0][0][5]~q ),
	.twiddle_data006(\twiddle_data[0][0][6]~q ),
	.twiddle_data007(\twiddle_data[0][0][7]~q ),
	.twiddle_data008(\twiddle_data[0][0][8]~q ),
	.twiddle_data009(\twiddle_data[0][0][9]~q ),
	.twiddle_data110(\twiddle_data[1][1][0]~q ),
	.twiddle_data111(\twiddle_data[1][1][1]~q ),
	.twiddle_data112(\twiddle_data[1][1][2]~q ),
	.twiddle_data113(\twiddle_data[1][1][3]~q ),
	.twiddle_data114(\twiddle_data[1][1][4]~q ),
	.twiddle_data115(\twiddle_data[1][1][5]~q ),
	.twiddle_data116(\twiddle_data[1][1][6]~q ),
	.twiddle_data117(\twiddle_data[1][1][7]~q ),
	.twiddle_data118(\twiddle_data[1][1][8]~q ),
	.twiddle_data119(\twiddle_data[1][1][9]~q ),
	.twiddle_data100(\twiddle_data[1][0][0]~q ),
	.twiddle_data101(\twiddle_data[1][0][1]~q ),
	.twiddle_data102(\twiddle_data[1][0][2]~q ),
	.twiddle_data103(\twiddle_data[1][0][3]~q ),
	.twiddle_data104(\twiddle_data[1][0][4]~q ),
	.twiddle_data105(\twiddle_data[1][0][5]~q ),
	.twiddle_data106(\twiddle_data[1][0][6]~q ),
	.twiddle_data107(\twiddle_data[1][0][7]~q ),
	.twiddle_data108(\twiddle_data[1][0][8]~q ),
	.twiddle_data109(\twiddle_data[1][0][9]~q ),
	.twiddle_data210(\twiddle_data[2][1][0]~q ),
	.twiddle_data211(\twiddle_data[2][1][1]~q ),
	.twiddle_data212(\twiddle_data[2][1][2]~q ),
	.twiddle_data213(\twiddle_data[2][1][3]~q ),
	.twiddle_data214(\twiddle_data[2][1][4]~q ),
	.twiddle_data215(\twiddle_data[2][1][5]~q ),
	.twiddle_data216(\twiddle_data[2][1][6]~q ),
	.twiddle_data217(\twiddle_data[2][1][7]~q ),
	.twiddle_data218(\twiddle_data[2][1][8]~q ),
	.twiddle_data219(\twiddle_data[2][1][9]~q ),
	.twiddle_data200(\twiddle_data[2][0][0]~q ),
	.twiddle_data201(\twiddle_data[2][0][1]~q ),
	.twiddle_data202(\twiddle_data[2][0][2]~q ),
	.twiddle_data203(\twiddle_data[2][0][3]~q ),
	.twiddle_data204(\twiddle_data[2][0][4]~q ),
	.twiddle_data205(\twiddle_data[2][0][5]~q ),
	.twiddle_data206(\twiddle_data[2][0][6]~q ),
	.twiddle_data207(\twiddle_data[2][0][7]~q ),
	.twiddle_data208(\twiddle_data[2][0][8]~q ),
	.twiddle_data209(\twiddle_data[2][0][9]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_cxb_data_r_1 ram_cxb_bfp_data(
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_8_0(\ram_cxb_bfp_data|ram_in_reg[0][8]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_8_2(\ram_cxb_bfp_data|ram_in_reg[2][8]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_8_1(\ram_cxb_bfp_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_8_3(\ram_cxb_bfp_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_9_0(\ram_cxb_bfp_data|ram_in_reg[0][9]~q ),
	.ram_in_reg_9_2(\ram_cxb_bfp_data|ram_in_reg[2][9]~q ),
	.ram_in_reg_9_1(\ram_cxb_bfp_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_3(\ram_cxb_bfp_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_8_4(\ram_cxb_bfp_data|ram_in_reg[4][8]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_8_6(\ram_cxb_bfp_data|ram_in_reg[6][8]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_8_5(\ram_cxb_bfp_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_8_7(\ram_cxb_bfp_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_9_4(\ram_cxb_bfp_data|ram_in_reg[4][9]~q ),
	.ram_in_reg_9_6(\ram_cxb_bfp_data|ram_in_reg[6][9]~q ),
	.ram_in_reg_9_5(\ram_cxb_bfp_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_9_7(\ram_cxb_bfp_data|ram_in_reg[7][9]~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.ram_data_out0_17(\ccc|ram_data_out0[17]~q ),
	.ram_data_out1_17(\ccc|ram_data_out1[17]~q ),
	.sw_r_tdl_0_4(\sw_r_tdl[4][0]~q ),
	.ram_data_out2_17(\ccc|ram_data_out2[17]~q ),
	.ram_data_out3_17(\ccc|ram_data_out3[17]~q ),
	.sw_r_tdl_1_4(\sw_r_tdl[4][1]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_16(\ccc|ram_data_out0[16]~q ),
	.ram_data_out1_16(\ccc|ram_data_out1[16]~q ),
	.ram_data_out2_16(\ccc|ram_data_out2[16]~q ),
	.ram_data_out3_16(\ccc|ram_data_out3[16]~q ),
	.ram_data_out0_18(\ccc|ram_data_out0[18]~q ),
	.ram_data_out1_18(\ccc|ram_data_out1[18]~q ),
	.ram_data_out2_18(\ccc|ram_data_out2[18]~q ),
	.ram_data_out3_18(\ccc|ram_data_out3[18]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.ram_data_out0_19(\ccc|ram_data_out0[19]~q ),
	.ram_data_out1_19(\ccc|ram_data_out1[19]~q ),
	.ram_data_out2_19(\ccc|ram_data_out2[19]~q ),
	.ram_data_out3_19(\ccc|ram_data_out3[19]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.clk(clk));

fftsign_asj_fft_cxb_data ram_cxb_wr_data(
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_9_3(\ram_cxb_wr_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_9_0(\ram_cxb_wr_data|ram_in_reg[0][9]~q ),
	.ram_in_reg_9_1(\ram_cxb_wr_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_2(\ram_cxb_wr_data|ram_in_reg[2][9]~q ),
	.ram_in_reg_9_7(\ram_cxb_wr_data|ram_in_reg[7][9]~q ),
	.ram_in_reg_9_4(\ram_cxb_wr_data|ram_in_reg[4][9]~q ),
	.ram_in_reg_9_5(\ram_cxb_wr_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_9_6(\ram_cxb_wr_data|ram_in_reg[6][9]~q ),
	.ram_in_reg_8_3(\ram_cxb_wr_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_8_0(\ram_cxb_wr_data|ram_in_reg[0][8]~q ),
	.ram_in_reg_8_1(\ram_cxb_wr_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_8_2(\ram_cxb_wr_data|ram_in_reg[2][8]~q ),
	.ram_in_reg_8_7(\ram_cxb_wr_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_8_4(\ram_cxb_wr_data|ram_in_reg[4][8]~q ),
	.ram_in_reg_8_5(\ram_cxb_wr_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_8_6(\ram_cxb_wr_data|ram_in_reg[6][8]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_block3a1(\get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_block3a0(\get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.reg_no_twiddle605(\bfpdft|reg_no_twiddle[6][0][5]~q ),
	.reg_no_twiddle609(\bfpdft|reg_no_twiddle[6][0][9]~q ),
	.reg_no_twiddle615(\bfpdft|reg_no_twiddle[6][1][5]~q ),
	.reg_no_twiddle619(\bfpdft|reg_no_twiddle[6][1][9]~q ),
	.tdl_arr_5_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][9]~q ),
	.tdl_arr_5_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_9_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][9]~q ),
	.reg_no_twiddle606(\bfpdft|reg_no_twiddle[6][0][6]~q ),
	.reg_no_twiddle616(\bfpdft|reg_no_twiddle[6][1][6]~q ),
	.tdl_arr_6_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][6]~q ),
	.reg_no_twiddle607(\bfpdft|reg_no_twiddle[6][0][7]~q ),
	.reg_no_twiddle617(\bfpdft|reg_no_twiddle[6][1][7]~q ),
	.tdl_arr_7_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_7_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][7]~q ),
	.reg_no_twiddle608(\bfpdft|reg_no_twiddle[6][0][8]~q ),
	.reg_no_twiddle618(\bfpdft|reg_no_twiddle[6][1][8]~q ),
	.tdl_arr_8_1(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_11(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_12(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_13(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_14(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][8]~q ),
	.tdl_arr_8_15(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][8]~q ),
	.tdl_arr_2_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][2]~q ),
	.reg_no_twiddle602(\bfpdft|reg_no_twiddle[6][0][2]~q ),
	.tdl_arr_2_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][2]~q ),
	.reg_no_twiddle612(\bfpdft|reg_no_twiddle[6][1][2]~q ),
	.tdl_arr_1_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][1]~q ),
	.reg_no_twiddle601(\bfpdft|reg_no_twiddle[6][0][1]~q ),
	.tdl_arr_1_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][1]~q ),
	.reg_no_twiddle611(\bfpdft|reg_no_twiddle[6][1][1]~q ),
	.tdl_arr_0_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][0]~q ),
	.reg_no_twiddle600(\bfpdft|reg_no_twiddle[6][0][0]~q ),
	.tdl_arr_0_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][0]~q ),
	.reg_no_twiddle610(\bfpdft|reg_no_twiddle[6][1][0]~q ),
	.tdl_arr_4_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][4]~q ),
	.reg_no_twiddle604(\bfpdft|reg_no_twiddle[6][0][4]~q ),
	.tdl_arr_4_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][4]~q ),
	.reg_no_twiddle614(\bfpdft|reg_no_twiddle[6][1][4]~q ),
	.tdl_arr_3_1(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_11(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_12(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:imag_delay|tdl_arr[1][3]~q ),
	.reg_no_twiddle603(\bfpdft|reg_no_twiddle[6][0][3]~q ),
	.tdl_arr_3_13(\bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_14(\bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_3_15(\bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:real_delay|tdl_arr[1][3]~q ),
	.reg_no_twiddle613(\bfpdft|reg_no_twiddle[6][1][3]~q ),
	.clk(clk));

fftsign_asj_fft_cxb_addr_2 ram_cxb_wr(
	.ram_in_reg_1_3(\ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr|ram_in_reg[3][5]~q ),
	.ram_block3a0(\ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a1(\ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_in_reg_1_0(\ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr|ram_in_reg[2][5]~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.ram_in_reg_0_1(\ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr|ram_in_reg[1][2]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr|ram_in_reg[1][4]~q ),
	.ram_in_reg_0_11(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_31(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_2_11(\ram_cxb_rd|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_31(\ram_cxb_rd|ram_in_reg[3][3]~q ),
	.ram_in_reg_4_11(\ram_cxb_rd|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_31(\ram_cxb_rd|ram_in_reg[3][5]~q ),
	.ram_in_reg_6_0(\ram_cxb_rd|ram_in_reg[0][6]~q ),
	.ram_in_reg_7_0(\ram_cxb_rd|ram_in_reg[0][7]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_0_01(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_01(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_01(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_01(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_01(\ram_cxb_rd|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_01(\ram_cxb_rd|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_11(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_3_11(\ram_cxb_rd|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_11(\ram_cxb_rd|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_21(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_21(\ram_cxb_rd|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_21(\ram_cxb_rd|ram_in_reg[2][5]~q ),
	.swa_tdl_0_16(\get_wr_swtiches|swa_tdl[16][0]~q ),
	.swa_tdl_1_16(\get_wr_swtiches|swa_tdl[16][1]~q ),
	.clk(clk));

fftsign_asj_fft_wrswgen get_wr_swtiches(
	.ram_block3a1(\get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_block3a0(\get_wr_swtiches|swd_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a2(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.ram_block3a3(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.swa_tdl_0_16(\get_wr_swtiches|swa_tdl[16][0]~q ),
	.swa_tdl_1_16(\get_wr_swtiches|swa_tdl[16][1]~q ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.Add1(\rd_adgen|Add1~0_combout ),
	.Mux1(\rd_adgen|Mux1~0_combout ),
	.Mux11(\rd_adgen|Mux1~1_combout ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.Add0(\rd_adgen|Add0~0_combout ),
	.Add11(\rd_adgen|Add1~1_combout ),
	.Add12(\rd_adgen|Add1~2_combout ),
	.Mux0(\rd_adgen|Mux0~0_combout ),
	.Mux01(\rd_adgen|Mux0~1_combout ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.clk(clk));

fftsign_asj_fft_cxb_addr_1 ram_cxb_rd(
	.global_clock_enable(\global_clock_enable~1_combout ),
	.ram_in_reg_0_1(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_2_1(\ram_cxb_rd|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_rd|ram_in_reg[3][3]~q ),
	.ram_in_reg_4_1(\ram_cxb_rd|ram_in_reg[1][4]~q ),
	.ram_in_reg_5_3(\ram_cxb_rd|ram_in_reg[3][5]~q ),
	.ram_in_reg_6_0(\ram_cxb_rd|ram_in_reg[0][6]~q ),
	.ram_in_reg_7_0(\ram_cxb_rd|ram_in_reg[0][7]~q ),
	.ram_in_reg_0_0(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\ram_cxb_rd|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_0(\ram_cxb_rd|ram_in_reg[0][5]~q ),
	.ram_in_reg_1_1(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_3_1(\ram_cxb_rd|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_1(\ram_cxb_rd|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_2(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_2(\ram_cxb_rd|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_rd|ram_in_reg[2][5]~q ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_c_2(\rd_adgen|rd_addr_c[2]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_b_3(\rd_adgen|rd_addr_b[3]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_c_4(\rd_adgen|rd_addr_c[4]~q ),
	.rd_addr_d_4(\rd_adgen|rd_addr_d[4]~q ),
	.rd_addr_b_5(\rd_adgen|rd_addr_b[5]~q ),
	.rd_addr_d_5(\rd_adgen|rd_addr_d[5]~q ),
	.rd_addr_d_6(\rd_adgen|rd_addr_d[6]~q ),
	.rd_addr_d_7(\rd_adgen|rd_addr_d[7]~q ),
	.clk(clk));

fftsign_asj_fft_dataadgen rd_adgen(
	.global_clock_enable(\global_clock_enable~1_combout ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_c_2(\rd_adgen|rd_addr_c[2]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_b_3(\rd_adgen|rd_addr_b[3]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_c_4(\rd_adgen|rd_addr_c[4]~q ),
	.rd_addr_d_4(\rd_adgen|rd_addr_d[4]~q ),
	.rd_addr_b_5(\rd_adgen|rd_addr_b[5]~q ),
	.rd_addr_d_5(\rd_adgen|rd_addr_d[5]~q ),
	.rd_addr_d_6(\rd_adgen|rd_addr_d[6]~q ),
	.rd_addr_d_7(\rd_adgen|rd_addr_d[7]~q ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.k_count_4(\ctrl|k_count[4]~q ),
	.k_count_0(\ctrl|k_count[0]~q ),
	.k_count_2(\ctrl|k_count[2]~q ),
	.Add1(\rd_adgen|Add1~0_combout ),
	.Mux1(\rd_adgen|Mux1~0_combout ),
	.Mux11(\rd_adgen|Mux1~1_combout ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.k_count_1(\ctrl|k_count[1]~q ),
	.k_count_3(\ctrl|k_count[3]~q ),
	.Add0(\rd_adgen|Add0~0_combout ),
	.k_count_5(\ctrl|k_count[5]~q ),
	.Add11(\rd_adgen|Add1~1_combout ),
	.Add12(\rd_adgen|Add1~2_combout ),
	.Mux0(\rd_adgen|Mux0~0_combout ),
	.Mux01(\rd_adgen|Mux0~1_combout ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.Mux02(\twid_factors|Mux0~0_combout ),
	.Mux12(\rd_adgen|Mux1~5_combout ),
	.Mux13(\rd_adgen|Mux1~6_combout ),
	.Mux03(\rd_adgen|Mux0~5_combout ),
	.Mux04(\rd_adgen|Mux0~6_combout ),
	.clk(clk));

fftsign_asj_fft_tdl_bit_2 \no_del_input_blk:delay_next_block (
	.data_in(\writer|rdy_for_next_block~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_0(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.clk(clk));

fftsign_asj_fft_tdl_bit_rst_6 delay_sop(
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_6(\delay_sop|tdl_arr[6]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_lpp_serial \gen_radix_4_last_pass:lpp (
	.ram_in_reg_2_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_1_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ),
	.data_3_imag_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][9]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][8]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q }),
	.data_1_imag_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][9]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][8]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q }),
	.ram_in_reg_9_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_9_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][9]~q ),
	.ram_in_reg_9_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_8_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_8_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_8_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_8_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_7_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_6_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_5_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_4_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_3_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ),
	.data_3_real_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][9]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][8]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q }),
	.data_1_real_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][9]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][8]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q }),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.data_imag_o_0(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.data_real_o_0(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.data_imag_o_1(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.data_real_o_1(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.data_imag_o_2(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.data_real_o_2(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.data_imag_o_3(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.data_real_o_3(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.data_imag_o_4(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.data_real_o_4(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.data_imag_o_5(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.data_real_o_5(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.data_imag_o_6(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.data_real_o_6(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.data_imag_o_7(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.data_real_o_7(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.data_imag_o_8(\gen_radix_4_last_pass:lpp|data_imag_o[8]~q ),
	.data_real_o_8(\gen_radix_4_last_pass:lpp|data_real_o[8]~q ),
	.data_imag_o_9(\gen_radix_4_last_pass:lpp|data_imag_o[9]~q ),
	.data_real_o_9(\gen_radix_4_last_pass:lpp|data_real_o[9]~q ),
	.wait_count_0(\sel_we|wait_count[0]~0_combout ),
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_41(\gen_radix_4_last_pass:lpp|gen_burst_val:delay_val|tdl_arr[4]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_cxb_data_r \gen_radix_4_last_pass:ram_cxb_lpp_data (
	.ram_in_reg_2_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_1_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_2_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_1_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_0_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_9_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_9_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][9]~q ),
	.ram_in_reg_9_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_8_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_8_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_8_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_8_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_7_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_6_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_5_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_4_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_3_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_9_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][9]~q ),
	.ram_in_reg_9_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][9]~q ),
	.ram_in_reg_8_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][8]~q ),
	.ram_in_reg_8_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][8]~q ),
	.ram_in_reg_7_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_6_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_5_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_4_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_3_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_2_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_1_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_9_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][9]~q ),
	.ram_in_reg_9_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][9]~q ),
	.ram_in_reg_8_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][8]~q ),
	.ram_in_reg_8_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][8]~q ),
	.ram_in_reg_7_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_6_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_5_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_4_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_3_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.lpp_ram_data_out_12_3(\lpp_ram_data_out[3][12]~q ),
	.lpp_ram_data_out_12_0(\lpp_ram_data_out[0][12]~q ),
	.tdl_arr_0_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.lpp_ram_data_out_12_1(\lpp_ram_data_out[1][12]~q ),
	.lpp_ram_data_out_12_2(\lpp_ram_data_out[2][12]~q ),
	.tdl_arr_1_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.lpp_ram_data_out_2_3(\lpp_ram_data_out[3][2]~q ),
	.lpp_ram_data_out_2_0(\lpp_ram_data_out[0][2]~q ),
	.lpp_ram_data_out_2_1(\lpp_ram_data_out[1][2]~q ),
	.lpp_ram_data_out_2_2(\lpp_ram_data_out[2][2]~q ),
	.lpp_ram_data_out_11_3(\lpp_ram_data_out[3][11]~q ),
	.lpp_ram_data_out_11_0(\lpp_ram_data_out[0][11]~q ),
	.lpp_ram_data_out_11_1(\lpp_ram_data_out[1][11]~q ),
	.lpp_ram_data_out_11_2(\lpp_ram_data_out[2][11]~q ),
	.lpp_ram_data_out_1_3(\lpp_ram_data_out[3][1]~q ),
	.lpp_ram_data_out_1_0(\lpp_ram_data_out[0][1]~q ),
	.lpp_ram_data_out_1_1(\lpp_ram_data_out[1][1]~q ),
	.lpp_ram_data_out_1_2(\lpp_ram_data_out[2][1]~q ),
	.lpp_ram_data_out_10_3(\lpp_ram_data_out[3][10]~q ),
	.lpp_ram_data_out_10_0(\lpp_ram_data_out[0][10]~q ),
	.lpp_ram_data_out_10_1(\lpp_ram_data_out[1][10]~q ),
	.lpp_ram_data_out_10_2(\lpp_ram_data_out[2][10]~q ),
	.lpp_ram_data_out_0_3(\lpp_ram_data_out[3][0]~q ),
	.lpp_ram_data_out_0_0(\lpp_ram_data_out[0][0]~q ),
	.lpp_ram_data_out_0_1(\lpp_ram_data_out[1][0]~q ),
	.lpp_ram_data_out_0_2(\lpp_ram_data_out[2][0]~q ),
	.lpp_ram_data_out_19_3(\lpp_ram_data_out[3][19]~q ),
	.lpp_ram_data_out_19_0(\lpp_ram_data_out[0][19]~q ),
	.lpp_ram_data_out_19_1(\lpp_ram_data_out[1][19]~q ),
	.lpp_ram_data_out_19_2(\lpp_ram_data_out[2][19]~q ),
	.lpp_ram_data_out_9_3(\lpp_ram_data_out[3][9]~q ),
	.lpp_ram_data_out_9_0(\lpp_ram_data_out[0][9]~q ),
	.lpp_ram_data_out_9_1(\lpp_ram_data_out[1][9]~q ),
	.lpp_ram_data_out_9_2(\lpp_ram_data_out[2][9]~q ),
	.lpp_ram_data_out_18_3(\lpp_ram_data_out[3][18]~q ),
	.lpp_ram_data_out_18_0(\lpp_ram_data_out[0][18]~q ),
	.lpp_ram_data_out_18_1(\lpp_ram_data_out[1][18]~q ),
	.lpp_ram_data_out_18_2(\lpp_ram_data_out[2][18]~q ),
	.lpp_ram_data_out_8_3(\lpp_ram_data_out[3][8]~q ),
	.lpp_ram_data_out_8_0(\lpp_ram_data_out[0][8]~q ),
	.lpp_ram_data_out_8_1(\lpp_ram_data_out[1][8]~q ),
	.lpp_ram_data_out_8_2(\lpp_ram_data_out[2][8]~q ),
	.lpp_ram_data_out_17_3(\lpp_ram_data_out[3][17]~q ),
	.lpp_ram_data_out_17_0(\lpp_ram_data_out[0][17]~q ),
	.lpp_ram_data_out_17_1(\lpp_ram_data_out[1][17]~q ),
	.lpp_ram_data_out_17_2(\lpp_ram_data_out[2][17]~q ),
	.lpp_ram_data_out_7_3(\lpp_ram_data_out[3][7]~q ),
	.lpp_ram_data_out_7_0(\lpp_ram_data_out[0][7]~q ),
	.lpp_ram_data_out_7_1(\lpp_ram_data_out[1][7]~q ),
	.lpp_ram_data_out_7_2(\lpp_ram_data_out[2][7]~q ),
	.lpp_ram_data_out_16_3(\lpp_ram_data_out[3][16]~q ),
	.lpp_ram_data_out_16_0(\lpp_ram_data_out[0][16]~q ),
	.lpp_ram_data_out_16_1(\lpp_ram_data_out[1][16]~q ),
	.lpp_ram_data_out_16_2(\lpp_ram_data_out[2][16]~q ),
	.lpp_ram_data_out_6_3(\lpp_ram_data_out[3][6]~q ),
	.lpp_ram_data_out_6_0(\lpp_ram_data_out[0][6]~q ),
	.lpp_ram_data_out_6_1(\lpp_ram_data_out[1][6]~q ),
	.lpp_ram_data_out_6_2(\lpp_ram_data_out[2][6]~q ),
	.lpp_ram_data_out_15_3(\lpp_ram_data_out[3][15]~q ),
	.lpp_ram_data_out_15_0(\lpp_ram_data_out[0][15]~q ),
	.lpp_ram_data_out_15_1(\lpp_ram_data_out[1][15]~q ),
	.lpp_ram_data_out_15_2(\lpp_ram_data_out[2][15]~q ),
	.lpp_ram_data_out_5_3(\lpp_ram_data_out[3][5]~q ),
	.lpp_ram_data_out_5_0(\lpp_ram_data_out[0][5]~q ),
	.lpp_ram_data_out_5_1(\lpp_ram_data_out[1][5]~q ),
	.lpp_ram_data_out_5_2(\lpp_ram_data_out[2][5]~q ),
	.lpp_ram_data_out_14_3(\lpp_ram_data_out[3][14]~q ),
	.lpp_ram_data_out_14_0(\lpp_ram_data_out[0][14]~q ),
	.lpp_ram_data_out_14_1(\lpp_ram_data_out[1][14]~q ),
	.lpp_ram_data_out_14_2(\lpp_ram_data_out[2][14]~q ),
	.lpp_ram_data_out_4_3(\lpp_ram_data_out[3][4]~q ),
	.lpp_ram_data_out_4_0(\lpp_ram_data_out[0][4]~q ),
	.lpp_ram_data_out_4_1(\lpp_ram_data_out[1][4]~q ),
	.lpp_ram_data_out_4_2(\lpp_ram_data_out[2][4]~q ),
	.lpp_ram_data_out_13_3(\lpp_ram_data_out[3][13]~q ),
	.lpp_ram_data_out_13_0(\lpp_ram_data_out[0][13]~q ),
	.lpp_ram_data_out_13_1(\lpp_ram_data_out[1][13]~q ),
	.lpp_ram_data_out_13_2(\lpp_ram_data_out[2][13]~q ),
	.lpp_ram_data_out_3_3(\lpp_ram_data_out[3][3]~q ),
	.lpp_ram_data_out_3_0(\lpp_ram_data_out[0][3]~q ),
	.lpp_ram_data_out_3_1(\lpp_ram_data_out[1][3]~q ),
	.lpp_ram_data_out_3_2(\lpp_ram_data_out[2][3]~q ),
	.clk(clk));

fftsign_asj_fft_cxb_addr \gen_radix_4_last_pass:ram_cxb_rd_lpp (
	.global_clock_enable(\global_clock_enable~1_combout ),
	.ram_in_reg_0_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_0(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ),
	.ram_in_reg_6_1(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ),
	.ram_in_reg_7_3(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_2(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[2][7]~q ),
	.rd_addr_d_0(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ),
	.rd_addr_d_1(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ),
	.rd_addr_d_2(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[2]~q ),
	.rd_addr_d_3(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[3]~q ),
	.rd_addr_d_4(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[4]~q ),
	.rd_addr_d_5(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[5]~q ),
	.sw_0(\gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ),
	.sw_1(\gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ),
	.clk(clk));

fftsign_asj_fft_lpprdadgen \gen_radix_4_last_pass:gen_lpp_addr (
	.lpp_c_i(\sel_we|lpp_c_i~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_0_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.tdl_arr_1_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.en_d1(\gen_radix_4_last_pass:gen_lpp_addr|en_d~q ),
	.rd_addr_d_0(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ),
	.rd_addr_d_1(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ),
	.rd_addr_d_2(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[2]~q ),
	.rd_addr_d_3(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[3]~q ),
	.rd_addr_d_4(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[4]~q ),
	.rd_addr_d_5(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[5]~q ),
	.sw_0(\gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ),
	.sw_1(\gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_3dp_rom twrom(
	.ram_block3a0(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a1(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.q_a_0(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_1(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_2(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_3(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_4(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_5(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_6(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_7(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_8(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_9(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.q_a_01(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_11(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_21(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_31(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_41(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_51(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_61(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_71(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_81(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_91(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.q_a_02(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_12(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_22(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_32(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_42(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_52(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_62(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_72(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_82(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_92(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.q_a_03(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_13(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_23(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_33(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_43(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_53(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_63(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_73(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_83(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_93(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.q_a_04(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_14(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_24(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_34(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_44(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_54(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_64(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_74(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_84(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_94(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.q_a_05(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_15(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_25(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_35(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_45(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_55(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_65(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_75(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_85(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.q_a_95(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.ram_block3a01(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a11(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_block3a2(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.ram_block3a3(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.ram_block3a4(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ),
	.ram_block3a5(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.clk(clk));

fftsign_asj_fft_twadgen twid_factors(
	.ram_block3a2(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.ram_block3a3(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.ram_block3a0(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a1(\twid_factors|twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_block3a01(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a11(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_block3a21(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.ram_block3a31(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.ram_block3a4(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ),
	.ram_block3a5(\twid_factors|twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.k_count_4(\ctrl|k_count[4]~q ),
	.k_count_2(\ctrl|k_count[2]~q ),
	.Mux1(\rd_adgen|Mux1~1_combout ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.k_count_3(\ctrl|k_count[3]~q ),
	.k_count_5(\ctrl|k_count[5]~q ),
	.Mux0(\rd_adgen|Mux0~1_combout ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.Mux01(\twid_factors|Mux0~0_combout ),
	.Mux11(\rd_adgen|Mux1~5_combout ),
	.Mux12(\rd_adgen|Mux1~6_combout ),
	.Mux02(\rd_adgen|Mux0~5_combout ),
	.Mux03(\rd_adgen|Mux0~6_combout ),
	.clk(clk));

fftsign_asj_fft_bfp_ctrl bfpc(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable1(\global_clock_enable~1_combout ),
	.blk_exp_0(\bfpc|blk_exp[0]~q ),
	.blk_exp_1(\bfpc|blk_exp[1]~q ),
	.blk_exp_2(\bfpc|blk_exp[2]~q ),
	.blk_exp_3(\bfpc|blk_exp[3]~q ),
	.blk_exp_4(\bfpc|blk_exp[4]~q ),
	.blk_exp_5(\bfpc|blk_exp[5]~q ),
	.exp_en(\exp_en~q ),
	.slb_last_0(\bfpc|slb_last[0]~q ),
	.slb_last_1(\bfpc|slb_last[1]~q ),
	.slb_last_2(\bfpc|slb_last[2]~q ),
	.slb_i_0(\bfpdft|gen_disc:bfp_detect|slb_i[0]~q ),
	.slb_i_1(\bfpdft|gen_disc:bfp_detect|slb_i[1]~q ),
	.slb_i_2(\bfpdft|gen_disc:bfp_detect|slb_i[2]~q ),
	.slb_i_3(\bfpdft|gen_disc:bfp_detect|slb_i[3]~q ),
	.Mux2(\bfpdft|gen_disc:bfp_detect|Mux2~0_combout ),
	.tdl_arr_23(\delay_blk_done|tdl_arr[23]~q ),
	.Mux1(\bfpdft|gen_disc:bfp_detect|Mux1~0_combout ),
	.tdl_arr_6(\bfpc|gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[6]~q ),
	.tdl_arr_9(\delay_np|tdl_arr[9]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_tdl_bit_3 delay_blk_done(
	.data_in(\ctrl|blk_done_int~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_23(\delay_blk_done|tdl_arr[23]~q ),
	.clk(clk));

fftsign_auk_dspip_avalon_streaming_sink auk_dsp_atlantic_sink_1(
	.q_b_2(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_12(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_1(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_11(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_0(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_10(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_9(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_19(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_8(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_18(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_7(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_17(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_6(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_16(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_5(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_15(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_4(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_14(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_3(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_13(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.at_sink_ready_s1(at_sink_ready_s),
	.send_eop_s1(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.sink_start1(\auk_dsp_atlantic_sink_1|sink_start~q ),
	.empty_dff(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_stall1(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.send_sop_s1(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.clk(clk),
	.reset_n(reset_n),
	.sink_valid(sink_valid),
	.sink_eop(sink_eop),
	.sink_sop(sink_sop),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.at_sink_data({sink_real[9],sink_real[8],sink_real[7],sink_real[6],sink_real[5],sink_real[4],sink_real[3],sink_real[2],sink_real[1],sink_real[0],sink_imag[9],sink_imag[8],sink_imag[7],sink_imag[6],sink_imag[5],sink_imag[4],sink_imag[3],sink_imag[2],sink_imag[1],sink_imag[0]}));

fftsign_asj_fft_4dp_ram dat_A(
	.q_b_12(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_2(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_11(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_1(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_13(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_14(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_15(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_10(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_0(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_19(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_191(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_192(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_193(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_9(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_18(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_181(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_182(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_183(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_8(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_17(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_171(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_172(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_173(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_7(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_16(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_161(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_162(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_163(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_6(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_151(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_154(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_5(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_141(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_144(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_4(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_131(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_134(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_3(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.wren_a_3(\wren_a[3]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_18(\ccc|wraddress_a_bus[18]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_20(\ccc|wraddress_a_bus[20]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.wraddress_a_bus_14(\ccc|wraddress_a_bus[14]~q ),
	.wraddress_a_bus_15(\ccc|wraddress_a_bus[15]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_18(\ccc|rdaddress_a_bus[18]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_20(\ccc|rdaddress_a_bus[20]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.rdaddress_a_bus_22(\ccc|rdaddress_a_bus[22]~q ),
	.rdaddress_a_bus_7(\ccc|rdaddress_a_bus[7]~q ),
	.wren_a_0(\wren_a[0]~q ),
	.a_ram_data_in_bus_72(\ccc|a_ram_data_in_bus[72]~q ),
	.wraddress_a_bus_24(\ccc|wraddress_a_bus[24]~q ),
	.wraddress_a_bus_25(\ccc|wraddress_a_bus[25]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_27(\ccc|wraddress_a_bus[27]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.wraddress_a_bus_29(\ccc|wraddress_a_bus[29]~q ),
	.rdaddress_a_bus_24(\ccc|rdaddress_a_bus[24]~q ),
	.rdaddress_a_bus_25(\ccc|rdaddress_a_bus[25]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_27(\ccc|rdaddress_a_bus[27]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.rdaddress_a_bus_29(\ccc|rdaddress_a_bus[29]~q ),
	.rdaddress_a_bus_14(\ccc|rdaddress_a_bus[14]~q ),
	.rdaddress_a_bus_31(\ccc|rdaddress_a_bus[31]~q ),
	.wren_a_1(\wren_a[1]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.wraddress_a_bus_17(\ccc|wraddress_a_bus[17]~q ),
	.wraddress_a_bus_19(\ccc|wraddress_a_bus[19]~q ),
	.wraddress_a_bus_21(\ccc|wraddress_a_bus[21]~q ),
	.rdaddress_a_bus_17(\ccc|rdaddress_a_bus[17]~q ),
	.rdaddress_a_bus_19(\ccc|rdaddress_a_bus[19]~q ),
	.rdaddress_a_bus_21(\ccc|rdaddress_a_bus[21]~q ),
	.rdaddress_a_bus_23(\ccc|rdaddress_a_bus[23]~q ),
	.wren_a_2(\wren_a[2]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.wraddress_a_bus_9(\ccc|wraddress_a_bus[9]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_9(\ccc|rdaddress_a_bus[9]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.rdaddress_a_bus_15(\ccc|rdaddress_a_bus[15]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_71(\ccc|a_ram_data_in_bus[71]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_70(\ccc|a_ram_data_in_bus[70]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_79(\ccc|a_ram_data_in_bus[79]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_69(\ccc|a_ram_data_in_bus[69]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_78(\ccc|a_ram_data_in_bus[78]~q ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_68(\ccc|a_ram_data_in_bus[68]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_77(\ccc|a_ram_data_in_bus[77]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_67(\ccc|a_ram_data_in_bus[67]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_76(\ccc|a_ram_data_in_bus[76]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_66(\ccc|a_ram_data_in_bus[66]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_75(\ccc|a_ram_data_in_bus[75]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_65(\ccc|a_ram_data_in_bus[65]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_74(\ccc|a_ram_data_in_bus[74]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_64(\ccc|a_ram_data_in_bus[64]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_73(\ccc|a_ram_data_in_bus[73]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.clk(clk));

fftsign_asj_fft_unbburst_ctrl ccc(
	.q_b_12(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_2(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_11(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_1(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_13(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_14(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_15(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_10(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_0(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_19(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_191(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_192(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_193(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.q_b_9(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_18(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_181(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_182(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_183(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.q_b_8(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_17(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_171(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_172(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_173(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.q_b_7(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_16(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_161(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_162(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_163(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.q_b_6(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_151(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_154(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_5(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_141(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_144(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_4(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_131(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_134(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_3(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.lpp_c_i(\sel_we|lpp_c_i~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr|ram_in_reg[3][3]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr|ram_in_reg[3][5]~q ),
	.ram_block3a0(\ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.ram_block3a1(\ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr|ram_in_reg[0][3]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr|ram_in_reg[0][5]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr|ram_in_reg[1][5]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr|ram_in_reg[2][5]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_1_31(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_01(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_11(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_21(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_9_3(\ram_cxb_wr_data|ram_in_reg[3][9]~q ),
	.ram_in_reg_9_0(\ram_cxb_wr_data|ram_in_reg[0][9]~q ),
	.ram_in_reg_9_1(\ram_cxb_wr_data|ram_in_reg[1][9]~q ),
	.ram_in_reg_9_2(\ram_cxb_wr_data|ram_in_reg[2][9]~q ),
	.ram_in_reg_9_7(\ram_cxb_wr_data|ram_in_reg[7][9]~q ),
	.ram_in_reg_9_4(\ram_cxb_wr_data|ram_in_reg[4][9]~q ),
	.ram_in_reg_9_5(\ram_cxb_wr_data|ram_in_reg[5][9]~q ),
	.ram_in_reg_9_6(\ram_cxb_wr_data|ram_in_reg[6][9]~q ),
	.ram_in_reg_8_3(\ram_cxb_wr_data|ram_in_reg[3][8]~q ),
	.ram_in_reg_8_0(\ram_cxb_wr_data|ram_in_reg[0][8]~q ),
	.ram_in_reg_8_1(\ram_cxb_wr_data|ram_in_reg[1][8]~q ),
	.ram_in_reg_8_2(\ram_cxb_wr_data|ram_in_reg[2][8]~q ),
	.ram_in_reg_8_7(\ram_cxb_wr_data|ram_in_reg[7][8]~q ),
	.ram_in_reg_8_4(\ram_cxb_wr_data|ram_in_reg[4][8]~q ),
	.ram_in_reg_8_5(\ram_cxb_wr_data|ram_in_reg[5][8]~q ),
	.ram_in_reg_8_6(\ram_cxb_wr_data|ram_in_reg[6][8]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_5_31(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_01(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_11(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_21(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_3_31(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_01(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_11(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_21(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.wraddress_a_bus_18(\ccc|wraddress_a_bus[18]~q ),
	.wraddress_a_bus_3(\ccc|wraddress_a_bus[3]~q ),
	.wraddress_a_bus_20(\ccc|wraddress_a_bus[20]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.wraddress_a_bus_14(\ccc|wraddress_a_bus[14]~q ),
	.wraddress_a_bus_15(\ccc|wraddress_a_bus[15]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.rdaddress_a_bus_18(\ccc|rdaddress_a_bus[18]~q ),
	.rdaddress_a_bus_3(\ccc|rdaddress_a_bus[3]~q ),
	.rdaddress_a_bus_20(\ccc|rdaddress_a_bus[20]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.rdaddress_a_bus_22(\ccc|rdaddress_a_bus[22]~q ),
	.rdaddress_a_bus_7(\ccc|rdaddress_a_bus[7]~q ),
	.a_ram_data_in_bus_72(\ccc|a_ram_data_in_bus[72]~q ),
	.wraddress_a_bus_24(\ccc|wraddress_a_bus[24]~q ),
	.wraddress_a_bus_25(\ccc|wraddress_a_bus[25]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_27(\ccc|wraddress_a_bus[27]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.wraddress_a_bus_29(\ccc|wraddress_a_bus[29]~q ),
	.rdaddress_a_bus_24(\ccc|rdaddress_a_bus[24]~q ),
	.rdaddress_a_bus_25(\ccc|rdaddress_a_bus[25]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_27(\ccc|rdaddress_a_bus[27]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.rdaddress_a_bus_29(\ccc|rdaddress_a_bus[29]~q ),
	.rdaddress_a_bus_14(\ccc|rdaddress_a_bus[14]~q ),
	.rdaddress_a_bus_31(\ccc|rdaddress_a_bus[31]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.wraddress_a_bus_17(\ccc|wraddress_a_bus[17]~q ),
	.wraddress_a_bus_19(\ccc|wraddress_a_bus[19]~q ),
	.wraddress_a_bus_21(\ccc|wraddress_a_bus[21]~q ),
	.rdaddress_a_bus_17(\ccc|rdaddress_a_bus[17]~q ),
	.rdaddress_a_bus_19(\ccc|rdaddress_a_bus[19]~q ),
	.rdaddress_a_bus_21(\ccc|rdaddress_a_bus[21]~q ),
	.rdaddress_a_bus_23(\ccc|rdaddress_a_bus[23]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.wraddress_a_bus_9(\ccc|wraddress_a_bus[9]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_9(\ccc|rdaddress_a_bus[9]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.rdaddress_a_bus_15(\ccc|rdaddress_a_bus[15]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_71(\ccc|a_ram_data_in_bus[71]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_70(\ccc|a_ram_data_in_bus[70]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_79(\ccc|a_ram_data_in_bus[79]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_69(\ccc|a_ram_data_in_bus[69]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_78(\ccc|a_ram_data_in_bus[78]~q ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_68(\ccc|a_ram_data_in_bus[68]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_77(\ccc|a_ram_data_in_bus[77]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_67(\ccc|a_ram_data_in_bus[67]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_76(\ccc|a_ram_data_in_bus[76]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_66(\ccc|a_ram_data_in_bus[66]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_75(\ccc|a_ram_data_in_bus[75]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_65(\ccc|a_ram_data_in_bus[65]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.a_ram_data_in_bus_74(\ccc|a_ram_data_in_bus[74]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_64(\ccc|a_ram_data_in_bus[64]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_73(\ccc|a_ram_data_in_bus[73]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.wc_vec_3(\wc_vec[3]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.sel_ram_in(\sel_ram_in~q ),
	.ram_in_reg_0_11(\ram_cxb_wr|ram_in_reg[1][0]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.data_rdy_vec_2(\data_rdy_vec[2]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.ram_in_reg_2_11(\ram_cxb_wr|ram_in_reg[1][2]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.ram_in_reg_4_11(\ram_cxb_wr|ram_in_reg[1][4]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.wr_address_i_int_7(\writer|wr_address_i_int[7]~q ),
	.ram_in_reg_0_12(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_01(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.data_rdy_vec_0(\data_rdy_vec[0]~q ),
	.ram_in_reg_1_32(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_02(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_12(\ram_cxb_rd|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_01(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_32(\ram_cxb_rd|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_02(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_12(\ram_cxb_rd|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_01(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_32(\ram_cxb_rd|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_02(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[0][5]~q ),
	.ram_in_reg_6_01(\ram_cxb_rd|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_11(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[1][6]~q ),
	.ram_in_reg_7_01(\ram_cxb_rd|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_31(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[3][7]~q ),
	.ram_in_reg_0_02(\ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_2_02(\ram_cxb_wr|ram_in_reg[0][2]~q ),
	.ram_in_reg_4_02(\ram_cxb_wr|ram_in_reg[0][4]~q ),
	.ram_in_reg_0_03(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_03(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_03(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_03(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_03(\ram_cxb_rd|ram_in_reg[0][4]~q ),
	.ram_in_reg_5_03(\ram_cxb_rd|ram_in_reg[0][5]~q ),
	.ram_in_reg_7_21(\gen_radix_4_last_pass:ram_cxb_rd_lpp|ram_in_reg[2][7]~q ),
	.ram_in_reg_1_12(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_3_12(\ram_cxb_rd|ram_in_reg[1][3]~q ),
	.ram_in_reg_5_12(\ram_cxb_rd|ram_in_reg[1][5]~q ),
	.ram_in_reg_1_22(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_3_22(\ram_cxb_rd|ram_in_reg[2][3]~q ),
	.ram_in_reg_5_22(\ram_cxb_rd|ram_in_reg[2][5]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.data_in_r_9(\writer|data_in_r[9]~q ),
	.data_in_i_9(\writer|data_in_i[9]~q ),
	.data_in_r_8(\writer|data_in_r[8]~q ),
	.data_in_i_8(\writer|data_in_i[8]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.ram_data_out0_17(\ccc|ram_data_out0[17]~q ),
	.ram_data_out1_17(\ccc|ram_data_out1[17]~q ),
	.ram_data_out2_17(\ccc|ram_data_out2[17]~q ),
	.ram_data_out3_17(\ccc|ram_data_out3[17]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_16(\ccc|ram_data_out0[16]~q ),
	.ram_data_out1_16(\ccc|ram_data_out1[16]~q ),
	.ram_data_out2_16(\ccc|ram_data_out2[16]~q ),
	.ram_data_out3_16(\ccc|ram_data_out3[16]~q ),
	.ram_data_out0_18(\ccc|ram_data_out0[18]~q ),
	.ram_data_out1_18(\ccc|ram_data_out1[18]~q ),
	.ram_data_out2_18(\ccc|ram_data_out2[18]~q ),
	.ram_data_out3_18(\ccc|ram_data_out3[18]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.ram_data_out0_19(\ccc|ram_data_out0[19]~q ),
	.ram_data_out1_19(\ccc|ram_data_out1[19]~q ),
	.ram_data_out2_19(\ccc|ram_data_out2[19]~q ),
	.ram_data_out3_19(\ccc|ram_data_out3[19]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.clk(clk));

fftsign_asj_fft_in_write_sgl writer(
	.rdy_for_next_block1(\writer|rdy_for_next_block~q ),
	.disable_wr1(\writer|disable_wr~q ),
	.data_rdy_int1(\writer|data_rdy_int~q ),
	.wren_3(\writer|wren[3]~q ),
	.wren_0(\writer|wren[0]~q ),
	.wren_1(\writer|wren[1]~q ),
	.wren_2(\writer|wren[2]~q ),
	.blk_done_int(\ctrl|blk_done_int~q ),
	.core_real_in_2(\core_real_in[2]~q ),
	.core_imag_in_2(\core_imag_in[2]~q ),
	.core_real_in_1(\core_real_in[1]~q ),
	.core_imag_in_1(\core_imag_in[1]~q ),
	.core_real_in_0(\core_real_in[0]~q ),
	.core_imag_in_0(\core_imag_in[0]~q ),
	.core_real_in_9(\core_real_in[9]~q ),
	.core_imag_in_9(\core_imag_in[9]~q ),
	.core_real_in_8(\core_real_in[8]~q ),
	.core_imag_in_8(\core_imag_in[8]~q ),
	.core_real_in_7(\core_real_in[7]~q ),
	.core_imag_in_7(\core_imag_in[7]~q ),
	.core_real_in_6(\core_real_in[6]~q ),
	.core_imag_in_6(\core_imag_in[6]~q ),
	.core_real_in_5(\core_real_in[5]~q ),
	.core_imag_in_5(\core_imag_in[5]~q ),
	.core_real_in_4(\core_real_in[4]~q ),
	.core_imag_in_4(\core_imag_in[4]~q ),
	.core_real_in_3(\core_real_in[3]~q ),
	.core_imag_in_3(\core_imag_in[3]~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wr_address_i_int_4(\writer|wr_address_i_int[4]~q ),
	.wr_address_i_int_5(\writer|wr_address_i_int[5]~q ),
	.wr_address_i_int_6(\writer|wr_address_i_int[6]~q ),
	.wr_address_i_int_7(\writer|wr_address_i_int[7]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.data_in_r_9(\writer|data_in_r[9]~q ),
	.data_in_i_9(\writer|data_in_i[9]~q ),
	.data_in_r_8(\writer|data_in_r[8]~q ),
	.data_in_i_8(\writer|data_in_i[8]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_wrengen sel_we(
	.lpp_c_i1(\sel_we|lpp_c_i~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.global_clock_enable1(\global_clock_enable~1_combout ),
	.wait_count_0(\sel_we|wait_count[0]~0_combout ),
	.wc_i_d1(\sel_we|wc_i_d~q ),
	.p_cd_en_2(\p_cd_en[2]~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_tdl_bit_rst_5 delay_np(
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_9(\delay_np|tdl_arr[9]~q ),
	.next_pass_i(\ctrl|next_pass_i~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_m_k_counter ctrl(
	.rdy_for_next_block(\writer|rdy_for_next_block~q ),
	.blk_done_int1(\ctrl|blk_done_int~q ),
	.global_clock_enable(\global_clock_enable~1_combout ),
	.tdl_arr_0(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.p_2(\ctrl|p[2]~q ),
	.p_0(\ctrl|p[0]~q ),
	.p_1(\ctrl|p[1]~q ),
	.k_count_4(\ctrl|k_count[4]~q ),
	.k_count_0(\ctrl|k_count[0]~q ),
	.k_count_2(\ctrl|k_count[2]~q ),
	.k_count_6(\ctrl|k_count[6]~q ),
	.k_count_1(\ctrl|k_count[1]~q ),
	.k_count_3(\ctrl|k_count[3]~q ),
	.k_count_5(\ctrl|k_count[5]~q ),
	.k_count_7(\ctrl|k_count[7]~q ),
	.data_rdy_vec_4(\data_rdy_vec[4]~q ),
	.next_pass_i1(\ctrl|next_pass_i~q ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_auk_dspip_avalon_streaming_controller auk_dsp_interface_controller_1(
	.master_sink_ena(\master_sink_ena~q ),
	.sink_in_work(\sink_in_work~q ),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_stall_reg1(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_stall_reg1(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.send_eop_s(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.sink_start(\auk_dsp_atlantic_sink_1|sink_start~q ),
	.empty_dff(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_stall(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.stall_reg1(\auk_dsp_interface_controller_1|stall_reg~q ),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

fftsign_auk_dspip_avalon_streaming_source auk_dsp_atlantic_source_1(
	.data_count({\data_count_sig[9]~q ,\data_count_sig[8]~q ,\data_count_sig[7]~q ,\data_count_sig[6]~q ,\data_count_sig[5]~q ,\data_count_sig[4]~q ,\data_count_sig[3]~q ,\data_count_sig[2]~q ,\data_count_sig[1]~q ,\data_count_sig[0]~q }),
	.at_source_valid_s1(at_source_valid_s),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s1(at_source_sop_s),
	.at_source_eop_s1(at_source_eop_s),
	.at_source_data_16(at_source_data_16),
	.at_source_data_17(at_source_data_17),
	.at_source_data_18(at_source_data_18),
	.at_source_data_19(at_source_data_19),
	.at_source_data_20(at_source_data_20),
	.at_source_data_21(at_source_data_21),
	.at_source_data_22(at_source_data_22),
	.at_source_data_23(at_source_data_23),
	.at_source_data_24(at_source_data_24),
	.at_source_data_25(at_source_data_25),
	.at_source_data_6(at_source_data_6),
	.at_source_data_7(at_source_data_7),
	.at_source_data_8(at_source_data_8),
	.at_source_data_9(at_source_data_9),
	.at_source_data_10(at_source_data_10),
	.at_source_data_11(at_source_data_11),
	.at_source_data_12(at_source_data_12),
	.at_source_data_13(at_source_data_13),
	.at_source_data_14(at_source_data_14),
	.at_source_data_15(at_source_data_15),
	.at_source_data_0(at_source_data_0),
	.at_source_data_1(at_source_data_1),
	.at_source_data_2(at_source_data_2),
	.at_source_data_3(at_source_data_3),
	.at_source_data_4(at_source_data_4),
	.at_source_data_5(at_source_data_5),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_stall_reg(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.master_source_ena(\master_source_ena~q ),
	.sink_ready_ctrl_d(\sink_ready_ctrl_d~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.sop(\sop~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.source_stall_int_d1(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.data({\fft_real_out[9]~q ,\fft_real_out[8]~q ,\fft_real_out[7]~q ,\fft_real_out[6]~q ,\fft_real_out[5]~q ,\fft_real_out[4]~q ,\fft_real_out[3]~q ,\fft_real_out[2]~q ,\fft_real_out[1]~q ,\fft_real_out[0]~q ,\fft_imag_out[9]~q ,\fft_imag_out[8]~q ,\fft_imag_out[7]~q ,
\fft_imag_out[6]~q ,\fft_imag_out[5]~q ,\fft_imag_out[4]~q ,\fft_imag_out[3]~q ,\fft_imag_out[2]~q ,\fft_imag_out[1]~q ,\fft_imag_out[0]~q ,\exponent_out[5]~q ,\exponent_out[4]~q ,\exponent_out[3]~q ,\exponent_out[2]~q ,\exponent_out[1]~q ,\exponent_out[0]~q }),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready));

dffeas master_sink_ena(
	.clk(clk),
	.d(\WideOr1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\master_sink_ena~q ),
	.prn(vcc));
defparam master_sink_ena.is_wysiwyg = "true";
defparam master_sink_ena.power_up = "low";

dffeas sink_in_work(
	.clk(clk),
	.d(\sink_in_work~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_in_work~q ),
	.prn(vcc));
defparam sink_in_work.is_wysiwyg = "true";
defparam sink_in_work.power_up = "low";

dffeas \data_count_sig[7] (
	.clk(clk),
	.d(\data_count_sig[7]~24_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[7]~q ),
	.prn(vcc));
defparam \data_count_sig[7] .is_wysiwyg = "true";
defparam \data_count_sig[7] .power_up = "low";

dffeas \data_count_sig[9] (
	.clk(clk),
	.d(\data_count_sig[9]~31_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[9]~q ),
	.prn(vcc));
defparam \data_count_sig[9] .is_wysiwyg = "true";
defparam \data_count_sig[9] .power_up = "low";

dffeas \data_count_sig[8] (
	.clk(clk),
	.d(\data_count_sig[8]~29_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[8]~q ),
	.prn(vcc));
defparam \data_count_sig[8] .is_wysiwyg = "true";
defparam \data_count_sig[8] .power_up = "low";

dffeas \data_count_sig[3] (
	.clk(clk),
	.d(\data_count_sig[3]~16_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[3]~q ),
	.prn(vcc));
defparam \data_count_sig[3] .is_wysiwyg = "true";
defparam \data_count_sig[3] .power_up = "low";

dffeas \data_count_sig[4] (
	.clk(clk),
	.d(\data_count_sig[4]~18_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[4]~q ),
	.prn(vcc));
defparam \data_count_sig[4] .is_wysiwyg = "true";
defparam \data_count_sig[4] .power_up = "low";

dffeas \data_count_sig[6] (
	.clk(clk),
	.d(\data_count_sig[6]~22_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[6]~q ),
	.prn(vcc));
defparam \data_count_sig[6] .is_wysiwyg = "true";
defparam \data_count_sig[6] .power_up = "low";

dffeas \data_count_sig[5] (
	.clk(clk),
	.d(\data_count_sig[5]~20_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[5]~q ),
	.prn(vcc));
defparam \data_count_sig[5] .is_wysiwyg = "true";
defparam \data_count_sig[5] .power_up = "low";

dffeas \data_count_sig[2] (
	.clk(clk),
	.d(\data_count_sig[2]~14_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[2]~q ),
	.prn(vcc));
defparam \data_count_sig[2] .is_wysiwyg = "true";
defparam \data_count_sig[2] .power_up = "low";

dffeas \data_count_sig[0] (
	.clk(clk),
	.d(\data_count_sig[0]~10_combout ),
	.asdata(\master_source_sop~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[0]~q ),
	.prn(vcc));
defparam \data_count_sig[0] .is_wysiwyg = "true";
defparam \data_count_sig[0] .power_up = "low";

dffeas \data_count_sig[1] (
	.clk(clk),
	.d(\data_count_sig[1]~12_combout ),
	.asdata(GND_port),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_count_sig[9]~27_combout ),
	.ena(\data_count_sig[3]~28_combout ),
	.q(\data_count_sig[1]~q ),
	.prn(vcc));
defparam \data_count_sig[1] .is_wysiwyg = "true";
defparam \data_count_sig[1] .power_up = "low";

cycloneive_lcell_comb \data_count_sig[0]~10 (
	.dataa(\data_count_sig[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\data_count_sig[0]~10_combout ),
	.cout(\data_count_sig[0]~11 ));
defparam \data_count_sig[0]~10 .lut_mask = 16'h55AA;
defparam \data_count_sig[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[1]~12 (
	.dataa(\data_count_sig[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[0]~11 ),
	.combout(\data_count_sig[1]~12_combout ),
	.cout(\data_count_sig[1]~13 ));
defparam \data_count_sig[1]~12 .lut_mask = 16'h5A5F;
defparam \data_count_sig[1]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[2]~14 (
	.dataa(\data_count_sig[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[1]~13 ),
	.combout(\data_count_sig[2]~14_combout ),
	.cout(\data_count_sig[2]~15 ));
defparam \data_count_sig[2]~14 .lut_mask = 16'h5AAF;
defparam \data_count_sig[2]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[3]~16 (
	.dataa(\data_count_sig[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[2]~15 ),
	.combout(\data_count_sig[3]~16_combout ),
	.cout(\data_count_sig[3]~17 ));
defparam \data_count_sig[3]~16 .lut_mask = 16'h5A5F;
defparam \data_count_sig[3]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[4]~18 (
	.dataa(\data_count_sig[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[3]~17 ),
	.combout(\data_count_sig[4]~18_combout ),
	.cout(\data_count_sig[4]~19 ));
defparam \data_count_sig[4]~18 .lut_mask = 16'h5AAF;
defparam \data_count_sig[4]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[5]~20 (
	.dataa(\data_count_sig[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[4]~19 ),
	.combout(\data_count_sig[5]~20_combout ),
	.cout(\data_count_sig[5]~21 ));
defparam \data_count_sig[5]~20 .lut_mask = 16'h5A5F;
defparam \data_count_sig[5]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[6]~22 (
	.dataa(\data_count_sig[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[5]~21 ),
	.combout(\data_count_sig[6]~22_combout ),
	.cout(\data_count_sig[6]~23 ));
defparam \data_count_sig[6]~22 .lut_mask = 16'h5AAF;
defparam \data_count_sig[6]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[7]~24 (
	.dataa(\data_count_sig[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[6]~23 ),
	.combout(\data_count_sig[7]~24_combout ),
	.cout(\data_count_sig[7]~25 ));
defparam \data_count_sig[7]~24 .lut_mask = 16'h5A5F;
defparam \data_count_sig[7]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[8]~29 (
	.dataa(\data_count_sig[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_count_sig[7]~25 ),
	.combout(\data_count_sig[8]~29_combout ),
	.cout(\data_count_sig[8]~30 ));
defparam \data_count_sig[8]~29 .lut_mask = 16'h5AAF;
defparam \data_count_sig[8]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_count_sig[9]~31 (
	.dataa(\data_count_sig[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\data_count_sig[8]~30 ),
	.combout(\data_count_sig[9]~31_combout ),
	.cout());
defparam \data_count_sig[9]~31 .lut_mask = 16'h5A5A;
defparam \data_count_sig[9]~31 .sum_lutc_input = "cin";

dffeas \core_real_in[2] (
	.clk(clk),
	.d(\core_real_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[2]~q ),
	.prn(vcc));
defparam \core_real_in[2] .is_wysiwyg = "true";
defparam \core_real_in[2] .power_up = "low";

dffeas \core_imag_in[2] (
	.clk(clk),
	.d(\core_imag_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[2]~q ),
	.prn(vcc));
defparam \core_imag_in[2] .is_wysiwyg = "true";
defparam \core_imag_in[2] .power_up = "low";

dffeas \core_real_in[1] (
	.clk(clk),
	.d(\core_real_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[1]~q ),
	.prn(vcc));
defparam \core_real_in[1] .is_wysiwyg = "true";
defparam \core_real_in[1] .power_up = "low";

dffeas \core_imag_in[1] (
	.clk(clk),
	.d(\core_imag_in~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[1]~q ),
	.prn(vcc));
defparam \core_imag_in[1] .is_wysiwyg = "true";
defparam \core_imag_in[1] .power_up = "low";

dffeas \core_real_in[0] (
	.clk(clk),
	.d(\core_real_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[0]~q ),
	.prn(vcc));
defparam \core_real_in[0] .is_wysiwyg = "true";
defparam \core_real_in[0] .power_up = "low";

dffeas \core_imag_in[0] (
	.clk(clk),
	.d(\core_imag_in~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[0]~q ),
	.prn(vcc));
defparam \core_imag_in[0] .is_wysiwyg = "true";
defparam \core_imag_in[0] .power_up = "low";

dffeas \core_real_in[9] (
	.clk(clk),
	.d(\core_real_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[9]~q ),
	.prn(vcc));
defparam \core_real_in[9] .is_wysiwyg = "true";
defparam \core_real_in[9] .power_up = "low";

dffeas \core_imag_in[9] (
	.clk(clk),
	.d(\core_imag_in~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[9]~q ),
	.prn(vcc));
defparam \core_imag_in[9] .is_wysiwyg = "true";
defparam \core_imag_in[9] .power_up = "low";

dffeas \core_real_in[8] (
	.clk(clk),
	.d(\core_real_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[8]~q ),
	.prn(vcc));
defparam \core_real_in[8] .is_wysiwyg = "true";
defparam \core_real_in[8] .power_up = "low";

dffeas \core_imag_in[8] (
	.clk(clk),
	.d(\core_imag_in~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[8]~q ),
	.prn(vcc));
defparam \core_imag_in[8] .is_wysiwyg = "true";
defparam \core_imag_in[8] .power_up = "low";

dffeas \core_real_in[7] (
	.clk(clk),
	.d(\core_real_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[7]~q ),
	.prn(vcc));
defparam \core_real_in[7] .is_wysiwyg = "true";
defparam \core_real_in[7] .power_up = "low";

dffeas \core_imag_in[7] (
	.clk(clk),
	.d(\core_imag_in~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[7]~q ),
	.prn(vcc));
defparam \core_imag_in[7] .is_wysiwyg = "true";
defparam \core_imag_in[7] .power_up = "low";

dffeas \core_real_in[6] (
	.clk(clk),
	.d(\core_real_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[6]~q ),
	.prn(vcc));
defparam \core_real_in[6] .is_wysiwyg = "true";
defparam \core_real_in[6] .power_up = "low";

dffeas \core_imag_in[6] (
	.clk(clk),
	.d(\core_imag_in~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[6]~q ),
	.prn(vcc));
defparam \core_imag_in[6] .is_wysiwyg = "true";
defparam \core_imag_in[6] .power_up = "low";

dffeas \core_real_in[5] (
	.clk(clk),
	.d(\core_real_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[5]~q ),
	.prn(vcc));
defparam \core_real_in[5] .is_wysiwyg = "true";
defparam \core_real_in[5] .power_up = "low";

dffeas \core_imag_in[5] (
	.clk(clk),
	.d(\core_imag_in~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[5]~q ),
	.prn(vcc));
defparam \core_imag_in[5] .is_wysiwyg = "true";
defparam \core_imag_in[5] .power_up = "low";

dffeas \core_real_in[4] (
	.clk(clk),
	.d(\core_real_in~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[4]~q ),
	.prn(vcc));
defparam \core_real_in[4] .is_wysiwyg = "true";
defparam \core_real_in[4] .power_up = "low";

dffeas \core_imag_in[4] (
	.clk(clk),
	.d(\core_imag_in~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[4]~q ),
	.prn(vcc));
defparam \core_imag_in[4] .is_wysiwyg = "true";
defparam \core_imag_in[4] .power_up = "low";

dffeas \core_real_in[3] (
	.clk(clk),
	.d(\core_real_in~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_real_in[3]~q ),
	.prn(vcc));
defparam \core_real_in[3] .is_wysiwyg = "true";
defparam \core_real_in[3] .power_up = "low";

dffeas \core_imag_in[3] (
	.clk(clk),
	.d(\core_imag_in~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\core_imag_in[3]~q ),
	.prn(vcc));
defparam \core_imag_in[3] .is_wysiwyg = "true";
defparam \core_imag_in[3] .power_up = "low";

dffeas master_source_ena(
	.clk(clk),
	.d(\master_source_ena~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\master_source_ena~q ),
	.prn(vcc));
defparam master_source_ena.is_wysiwyg = "true";
defparam master_source_ena.power_up = "low";

dffeas sink_ready_ctrl_d(
	.clk(clk),
	.d(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_ready_ctrl_d~q ),
	.prn(vcc));
defparam sink_ready_ctrl_d.is_wysiwyg = "true";
defparam sink_ready_ctrl_d.power_up = "low";

dffeas sop(
	.clk(clk),
	.d(\sop~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sop~q ),
	.prn(vcc));
defparam sop.is_wysiwyg = "true";
defparam sop.power_up = "low";

cycloneive_lcell_comb \global_clock_enable~0 (
	.dataa(gnd),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\global_clock_enable~0_combout ),
	.cout());
defparam \global_clock_enable~0 .lut_mask = 16'h3FFF;
defparam \global_clock_enable~0 .sum_lutc_input = "datac";

dffeas \fft_real_out[0] (
	.clk(clk),
	.d(\fft_real_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[0]~q ),
	.prn(vcc));
defparam \fft_real_out[0] .is_wysiwyg = "true";
defparam \fft_real_out[0] .power_up = "low";

dffeas \fft_real_out[1] (
	.clk(clk),
	.d(\fft_real_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[1]~q ),
	.prn(vcc));
defparam \fft_real_out[1] .is_wysiwyg = "true";
defparam \fft_real_out[1] .power_up = "low";

dffeas \fft_real_out[2] (
	.clk(clk),
	.d(\fft_real_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[2]~q ),
	.prn(vcc));
defparam \fft_real_out[2] .is_wysiwyg = "true";
defparam \fft_real_out[2] .power_up = "low";

dffeas \fft_real_out[3] (
	.clk(clk),
	.d(\fft_real_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[3]~q ),
	.prn(vcc));
defparam \fft_real_out[3] .is_wysiwyg = "true";
defparam \fft_real_out[3] .power_up = "low";

dffeas \fft_real_out[4] (
	.clk(clk),
	.d(\fft_real_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[4]~q ),
	.prn(vcc));
defparam \fft_real_out[4] .is_wysiwyg = "true";
defparam \fft_real_out[4] .power_up = "low";

dffeas \fft_real_out[5] (
	.clk(clk),
	.d(\fft_real_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[5]~q ),
	.prn(vcc));
defparam \fft_real_out[5] .is_wysiwyg = "true";
defparam \fft_real_out[5] .power_up = "low";

dffeas \fft_real_out[6] (
	.clk(clk),
	.d(\fft_real_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[6]~q ),
	.prn(vcc));
defparam \fft_real_out[6] .is_wysiwyg = "true";
defparam \fft_real_out[6] .power_up = "low";

dffeas \fft_real_out[7] (
	.clk(clk),
	.d(\fft_real_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[7]~q ),
	.prn(vcc));
defparam \fft_real_out[7] .is_wysiwyg = "true";
defparam \fft_real_out[7] .power_up = "low";

dffeas \fft_real_out[8] (
	.clk(clk),
	.d(\fft_real_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[8]~q ),
	.prn(vcc));
defparam \fft_real_out[8] .is_wysiwyg = "true";
defparam \fft_real_out[8] .power_up = "low";

dffeas \fft_real_out[9] (
	.clk(clk),
	.d(\fft_real_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_real_out[9]~q ),
	.prn(vcc));
defparam \fft_real_out[9] .is_wysiwyg = "true";
defparam \fft_real_out[9] .power_up = "low";

dffeas \fft_imag_out[0] (
	.clk(clk),
	.d(\fft_imag_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[0]~q ),
	.prn(vcc));
defparam \fft_imag_out[0] .is_wysiwyg = "true";
defparam \fft_imag_out[0] .power_up = "low";

dffeas \fft_imag_out[1] (
	.clk(clk),
	.d(\fft_imag_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[1]~q ),
	.prn(vcc));
defparam \fft_imag_out[1] .is_wysiwyg = "true";
defparam \fft_imag_out[1] .power_up = "low";

dffeas \fft_imag_out[2] (
	.clk(clk),
	.d(\fft_imag_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[2]~q ),
	.prn(vcc));
defparam \fft_imag_out[2] .is_wysiwyg = "true";
defparam \fft_imag_out[2] .power_up = "low";

dffeas \fft_imag_out[3] (
	.clk(clk),
	.d(\fft_imag_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[3]~q ),
	.prn(vcc));
defparam \fft_imag_out[3] .is_wysiwyg = "true";
defparam \fft_imag_out[3] .power_up = "low";

dffeas \fft_imag_out[4] (
	.clk(clk),
	.d(\fft_imag_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[4]~q ),
	.prn(vcc));
defparam \fft_imag_out[4] .is_wysiwyg = "true";
defparam \fft_imag_out[4] .power_up = "low";

dffeas \fft_imag_out[5] (
	.clk(clk),
	.d(\fft_imag_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[5]~q ),
	.prn(vcc));
defparam \fft_imag_out[5] .is_wysiwyg = "true";
defparam \fft_imag_out[5] .power_up = "low";

dffeas \fft_imag_out[6] (
	.clk(clk),
	.d(\fft_imag_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[6]~q ),
	.prn(vcc));
defparam \fft_imag_out[6] .is_wysiwyg = "true";
defparam \fft_imag_out[6] .power_up = "low";

dffeas \fft_imag_out[7] (
	.clk(clk),
	.d(\fft_imag_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[7]~q ),
	.prn(vcc));
defparam \fft_imag_out[7] .is_wysiwyg = "true";
defparam \fft_imag_out[7] .power_up = "low";

dffeas \fft_imag_out[8] (
	.clk(clk),
	.d(\fft_imag_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[8]~q ),
	.prn(vcc));
defparam \fft_imag_out[8] .is_wysiwyg = "true";
defparam \fft_imag_out[8] .power_up = "low";

dffeas \fft_imag_out[9] (
	.clk(clk),
	.d(\fft_imag_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_imag_out[9]~q ),
	.prn(vcc));
defparam \fft_imag_out[9] .is_wysiwyg = "true";
defparam \fft_imag_out[9] .power_up = "low";

dffeas \exponent_out[0] (
	.clk(clk),
	.d(\exponent_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[0]~q ),
	.prn(vcc));
defparam \exponent_out[0] .is_wysiwyg = "true";
defparam \exponent_out[0] .power_up = "low";

dffeas \exponent_out[1] (
	.clk(clk),
	.d(\exponent_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[1]~q ),
	.prn(vcc));
defparam \exponent_out[1] .is_wysiwyg = "true";
defparam \exponent_out[1] .power_up = "low";

dffeas \exponent_out[2] (
	.clk(clk),
	.d(\exponent_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[2]~q ),
	.prn(vcc));
defparam \exponent_out[2] .is_wysiwyg = "true";
defparam \exponent_out[2] .power_up = "low";

dffeas \exponent_out[3] (
	.clk(clk),
	.d(\exponent_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[3]~q ),
	.prn(vcc));
defparam \exponent_out[3] .is_wysiwyg = "true";
defparam \exponent_out[3] .power_up = "low";

dffeas \exponent_out[4] (
	.clk(clk),
	.d(\exponent_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[4]~q ),
	.prn(vcc));
defparam \exponent_out[4] .is_wysiwyg = "true";
defparam \exponent_out[4] .power_up = "low";

dffeas \exponent_out[5] (
	.clk(clk),
	.d(\exponent_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exponent_out[5]~q ),
	.prn(vcc));
defparam \exponent_out[5] .is_wysiwyg = "true";
defparam \exponent_out[5] .power_up = "low";

dffeas \fft_s1_cur.WAIT_FOR_INPUT (
	.clk(clk),
	.d(\fft_s1_cur.WAIT_FOR_INPUT~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.prn(vcc));
defparam \fft_s1_cur.WAIT_FOR_INPUT .is_wysiwyg = "true";
defparam \fft_s1_cur.WAIT_FOR_INPUT .power_up = "low";

dffeas \fft_s1_cur.WRITE_INPUT (
	.clk(clk),
	.d(\fft_s1_cur.WRITE_INPUT~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.WRITE_INPUT~q ),
	.prn(vcc));
defparam \fft_s1_cur.WRITE_INPUT .is_wysiwyg = "true";
defparam \fft_s1_cur.WRITE_INPUT .power_up = "low";

dffeas \fft_s1_cur.IDLE (
	.clk(clk),
	.d(\fft_s1_cur.WAIT_FOR_INPUT~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.IDLE~q ),
	.prn(vcc));
defparam \fft_s1_cur.IDLE .is_wysiwyg = "true";
defparam \fft_s1_cur.IDLE .power_up = "low";

cycloneive_lcell_comb \WideOr1~0 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(gnd),
	.datad(\fft_s1_cur.IDLE~q ),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hEEFF;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \global_clock_enable~1 (
	.dataa(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datab(\global_clock_enable~0_combout ),
	.datac(gnd),
	.datad(\auk_dsp_interface_controller_1|stall_reg~q ),
	.cin(gnd),
	.combout(\global_clock_enable~1_combout ),
	.cout());
defparam \global_clock_enable~1 .lut_mask = 16'hDD11;
defparam \global_clock_enable~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_in_work~0 (
	.dataa(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datab(\sink_in_work~q ),
	.datac(gnd),
	.datad(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.cin(gnd),
	.combout(\sink_in_work~0_combout ),
	.cout());
defparam \sink_in_work~0 .lut_mask = 16'hEEFF;
defparam \sink_in_work~0 .sum_lutc_input = "datac";

dffeas val_out(
	.clk(clk),
	.d(\val_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\val_out~q ),
	.prn(vcc));
defparam val_out.is_wysiwyg = "true";
defparam val_out.power_up = "low";

dffeas oe(
	.clk(clk),
	.d(\val_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\oe~q ),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

cycloneive_lcell_comb \master_source_ena~0 (
	.dataa(reset_n),
	.datab(\val_out~q ),
	.datac(\oe~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_ena~0_combout ),
	.cout());
defparam \master_source_ena~0 .lut_mask = 16'hFEFE;
defparam \master_source_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop~0 (
	.dataa(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.datab(\sink_ready_ctrl_d~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\sop~q ),
	.cin(gnd),
	.combout(\sop~0_combout ),
	.cout());
defparam \sop~0 .lut_mask = 16'hF7D5;
defparam \sop~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(\data_count_sig[3]~q ),
	.datab(\data_count_sig[9]~q ),
	.datac(\data_count_sig[8]~q ),
	.datad(\data_count_sig[7]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\data_count_sig[6]~q ),
	.datab(\data_count_sig[5]~q ),
	.datac(\data_count_sig[4]~q ),
	.datad(\data_count_sig[2]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\data_count_sig[1]~q ),
	.datad(\data_count_sig[0]~q ),
	.cin(gnd),
	.combout(\LessThan0~2_combout ),
	.cout());
defparam \LessThan0~2 .lut_mask = 16'h0FFF;
defparam \LessThan0~2 .sum_lutc_input = "datac";

dffeas master_source_sop(
	.clk(clk),
	.d(\master_source_sop~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\master_source_sop~q ),
	.prn(vcc));
defparam master_source_sop.is_wysiwyg = "true";
defparam master_source_sop.power_up = "low";

cycloneive_lcell_comb \data_count_sig[9]~26 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(\LessThan0~2_combout ),
	.datad(\master_source_sop~q ),
	.cin(gnd),
	.combout(\data_count_sig[9]~26_combout ),
	.cout());
defparam \data_count_sig[9]~26 .lut_mask = 16'hFEFF;
defparam \data_count_sig[9]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\data_count_sig[3]~q ),
	.datab(\data_count_sig[9]~q ),
	.datac(\data_count_sig[8]~q ),
	.datad(\data_count_sig[7]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\data_count_sig[6]~q ),
	.datab(\data_count_sig[5]~q ),
	.datac(\data_count_sig[4]~q ),
	.datad(\data_count_sig[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\data_count_sig[1]~q ),
	.datad(\data_count_sig[0]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[9]~27 (
	.dataa(\data_count_sig[9]~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\data_count_sig[9]~27_combout ),
	.cout());
defparam \data_count_sig[9]~27 .lut_mask = 16'hFF55;
defparam \data_count_sig[9]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_count_sig[3]~28 (
	.dataa(\global_clock_enable~1_combout ),
	.datab(\data_count_sig[9]~26_combout ),
	.datac(\Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_count_sig[3]~28_combout ),
	.cout());
defparam \data_count_sig[3]~28 .lut_mask = 16'hBFBF;
defparam \data_count_sig[3]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out[2]~0 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out[2]~0_combout ),
	.cout());
defparam \exponent_out[2]~0 .lut_mask = 16'hEEEE;
defparam \exponent_out[2]~0 .sum_lutc_input = "datac";

dffeas fft_dirn(
	.clk(clk),
	.d(\fft_dirn~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fft_dirn~q ),
	.prn(vcc));
defparam fft_dirn.is_wysiwyg = "true";
defparam fft_dirn.power_up = "low";

cycloneive_lcell_comb \fft_real_out~0 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~0_combout ),
	.cout());
defparam \fft_real_out~0 .lut_mask = 16'hFAFC;
defparam \fft_real_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~1 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~1_combout ),
	.cout());
defparam \fft_real_out~1 .lut_mask = 16'hFAFC;
defparam \fft_real_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~2 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~2_combout ),
	.cout());
defparam \fft_real_out~2 .lut_mask = 16'hFAFC;
defparam \fft_real_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~3 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~3_combout ),
	.cout());
defparam \fft_real_out~3 .lut_mask = 16'hFAFC;
defparam \fft_real_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~4 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~4_combout ),
	.cout());
defparam \fft_real_out~4 .lut_mask = 16'hFAFC;
defparam \fft_real_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~5 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~5_combout ),
	.cout());
defparam \fft_real_out~5 .lut_mask = 16'hFAFC;
defparam \fft_real_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~6 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~6_combout ),
	.cout());
defparam \fft_real_out~6 .lut_mask = 16'hFAFC;
defparam \fft_real_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~7 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~7_combout ),
	.cout());
defparam \fft_real_out~7 .lut_mask = 16'hFAFC;
defparam \fft_real_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~8 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[8]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[8]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~8_combout ),
	.cout());
defparam \fft_real_out~8 .lut_mask = 16'hFAFC;
defparam \fft_real_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_real_out~9 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_imag_o[9]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_real_o[9]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_real_out~9_combout ),
	.cout());
defparam \fft_real_out~9 .lut_mask = 16'hFAFC;
defparam \fft_real_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~0 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~0_combout ),
	.cout());
defparam \fft_imag_out~0 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~1 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~1_combout ),
	.cout());
defparam \fft_imag_out~1 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~2 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~2_combout ),
	.cout());
defparam \fft_imag_out~2 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~3 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~3_combout ),
	.cout());
defparam \fft_imag_out~3 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~4 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~4_combout ),
	.cout());
defparam \fft_imag_out~4 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~5 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~5_combout ),
	.cout());
defparam \fft_imag_out~5 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~6 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~6_combout ),
	.cout());
defparam \fft_imag_out~6 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~7 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~7_combout ),
	.cout());
defparam \fft_imag_out~7 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~8 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[8]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[8]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~8_combout ),
	.cout());
defparam \fft_imag_out~8 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_imag_out~9 (
	.dataa(\exponent_out[2]~0_combout ),
	.datab(\gen_radix_4_last_pass:lpp|data_real_o[9]~q ),
	.datac(\gen_radix_4_last_pass:lpp|data_imag_o[9]~q ),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\fft_imag_out~9_combout ),
	.cout());
defparam \fft_imag_out~9 .lut_mask = 16'hFAFC;
defparam \fft_imag_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~1 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~1_combout ),
	.cout());
defparam \exponent_out~1 .lut_mask = 16'hFEFE;
defparam \exponent_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~2 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~2_combout ),
	.cout());
defparam \exponent_out~2 .lut_mask = 16'hFEFE;
defparam \exponent_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~3 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~3_combout ),
	.cout());
defparam \exponent_out~3 .lut_mask = 16'hFEFE;
defparam \exponent_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~4 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~4_combout ),
	.cout());
defparam \exponent_out~4 .lut_mask = 16'hFEFE;
defparam \exponent_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~5 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~5_combout ),
	.cout());
defparam \exponent_out~5 .lut_mask = 16'hFEFE;
defparam \exponent_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \exponent_out~6 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\bfpc|blk_exp[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\exponent_out~6_combout ),
	.cout());
defparam \exponent_out~6 .lut_mask = 16'hFEFE;
defparam \exponent_out~6 .sum_lutc_input = "datac";

dffeas \fft_s1_cur.NO_WRITE (
	.clk(clk),
	.d(\fft_s1_cur.NO_WRITE~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.NO_WRITE~q ),
	.prn(vcc));
defparam \fft_s1_cur.NO_WRITE .is_wysiwyg = "true";
defparam \fft_s1_cur.NO_WRITE .power_up = "low";

dffeas \fft_s1_cur.DONE_WRITING (
	.clk(clk),
	.d(\fft_s1_cur.DONE_WRITING~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.DONE_WRITING~q ),
	.prn(vcc));
defparam \fft_s1_cur.DONE_WRITING .is_wysiwyg = "true";
defparam \fft_s1_cur.DONE_WRITING .power_up = "low";

dffeas \fft_s1_cur.EARLY_DONE (
	.clk(clk),
	.d(\fft_s1_cur.EARLY_DONE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.EARLY_DONE~q ),
	.prn(vcc));
defparam \fft_s1_cur.EARLY_DONE .is_wysiwyg = "true";
defparam \fft_s1_cur.EARLY_DONE .power_up = "low";

cycloneive_lcell_comb \fft_s1_cur.WAIT_FOR_INPUT~0 (
	.dataa(\fft_s1_cur.WRITE_INPUT~q ),
	.datab(\fft_s1_cur.NO_WRITE~q ),
	.datac(\fft_s1_cur.DONE_WRITING~q ),
	.datad(\fft_s1_cur.EARLY_DONE~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.WAIT_FOR_INPUT~0_combout ),
	.cout());
defparam \fft_s1_cur.WAIT_FOR_INPUT~0 .lut_mask = 16'h7FFF;
defparam \fft_s1_cur.WAIT_FOR_INPUT~0 .sum_lutc_input = "datac";

dffeas \fft_s1_cur.FFT_PROCESS_A (
	.clk(clk),
	.d(\fft_s1_cur.FFT_PROCESS_A~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s1_cur.NO_WRITE~4_combout ),
	.q(\fft_s1_cur.FFT_PROCESS_A~q ),
	.prn(vcc));
defparam \fft_s1_cur.FFT_PROCESS_A .is_wysiwyg = "true";
defparam \fft_s1_cur.FFT_PROCESS_A .power_up = "low";

cycloneive_lcell_comb \fft_s1_cur.WAIT_FOR_INPUT~1 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.WAIT_FOR_INPUT~0_combout ),
	.datac(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datad(\fft_s1_cur.FFT_PROCESS_A~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.WAIT_FOR_INPUT~1_combout ),
	.cout());
defparam \fft_s1_cur.WAIT_FOR_INPUT~1 .lut_mask = 16'hEFFF;
defparam \fft_s1_cur.WAIT_FOR_INPUT~1 .sum_lutc_input = "datac";

dffeas eop_out(
	.clk(clk),
	.d(\eop_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\eop_out~q ),
	.prn(vcc));
defparam eop_out.is_wysiwyg = "true";
defparam eop_out.power_up = "low";

dffeas \data_rdy_vec[24] (
	.clk(clk),
	.d(\data_rdy_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[24]~q ),
	.prn(vcc));
defparam \data_rdy_vec[24] .is_wysiwyg = "true";
defparam \data_rdy_vec[24] .power_up = "low";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~0 (
	.dataa(\fft_s1_cur.FFT_PROCESS_A~q ),
	.datab(\fft_s1_cur.NO_WRITE~q ),
	.datac(\eop_out~q ),
	.datad(\data_rdy_vec[24]~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~0_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~0 .lut_mask = 16'hEFFF;
defparam \fft_s1_cur.NO_WRITE~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~1 (
	.dataa(\fft_s1_cur.DONE_WRITING~q ),
	.datab(\fft_s1_cur.EARLY_DONE~q ),
	.datac(\no_del_input_blk:delay_next_block|tdl_arr[0]~q ),
	.datad(\writer|rdy_for_next_block~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~1_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~1 .lut_mask = 16'hEFFF;
defparam \fft_s1_cur.NO_WRITE~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~2 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\writer|disable_wr~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~2_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~2 .lut_mask = 16'hEFFF;
defparam \fft_s1_cur.NO_WRITE~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~3 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.NO_WRITE~0_combout ),
	.datac(\fft_s1_cur.NO_WRITE~1_combout ),
	.datad(\fft_s1_cur.NO_WRITE~2_combout ),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~3_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~3 .lut_mask = 16'hFFFE;
defparam \fft_s1_cur.NO_WRITE~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.WAIT_FOR_INPUT~2 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datab(\fft_s1_cur.WAIT_FOR_INPUT~1_combout ),
	.datac(\global_clock_enable~1_combout ),
	.datad(\fft_s1_cur.NO_WRITE~3_combout ),
	.cin(gnd),
	.combout(\fft_s1_cur.WAIT_FOR_INPUT~2_combout ),
	.cout());
defparam \fft_s1_cur.WAIT_FOR_INPUT~2 .lut_mask = 16'hEFFE;
defparam \fft_s1_cur.WAIT_FOR_INPUT~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.WRITE_INPUT~0 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.WAIT_FOR_INPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s1_cur.WRITE_INPUT~0_combout ),
	.cout());
defparam \fft_s1_cur.WRITE_INPUT~0 .lut_mask = 16'hEEEE;
defparam \fft_s1_cur.WRITE_INPUT~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~4 (
	.dataa(\fft_s1_cur.NO_WRITE~3_combout ),
	.datab(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datac(\global_clock_enable~0_combout ),
	.datad(\auk_dsp_interface_controller_1|stall_reg~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~4_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~4 .lut_mask = 16'hF737;
defparam \fft_s1_cur.NO_WRITE~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.WAIT_FOR_INPUT~3 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\fft_s1_cur.FFT_PROCESS_A~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.WAIT_FOR_INPUT~3_combout ),
	.cout());
defparam \fft_s1_cur.WAIT_FOR_INPUT~3 .lut_mask = 16'hAAFF;
defparam \fft_s1_cur.WAIT_FOR_INPUT~3 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.START_LPP (
	.clk(clk),
	.d(\fft_s2_cur.START_LPP~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.WAIT_FOR_LPP_INPUT~1_combout ),
	.q(\fft_s2_cur.START_LPP~q ),
	.prn(vcc));
defparam \fft_s2_cur.START_LPP .is_wysiwyg = "true";
defparam \fft_s2_cur.START_LPP .power_up = "low";

dffeas \fft_s2_cur.WAIT_FOR_LPP_INPUT (
	.clk(clk),
	.d(\fft_s2_cur.WAIT_FOR_LPP_INPUT~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.WAIT_FOR_LPP_INPUT~1_combout ),
	.q(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .power_up = "low";

cycloneive_lcell_comb \val_out~0 (
	.dataa(\fft_s2_cur.START_LPP~q ),
	.datab(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(gnd),
	.datad(\bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ),
	.cin(gnd),
	.combout(\val_out~0_combout ),
	.cout());
defparam \val_out~0 .lut_mask = 16'hFF77;
defparam \val_out~0 .sum_lutc_input = "datac";

dffeas \fft_s2_cur.LPP_OUTPUT_RDY (
	.clk(clk),
	.d(\fft_s2_cur.LPP_OUTPUT_RDY~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_OUTPUT_RDY .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_OUTPUT_RDY .power_up = "low";

dffeas \fft_s2_cur.LPP_DONE (
	.clk(clk),
	.d(\fft_s2_cur.LPP_DONE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\fft_s2_cur.LPP_DONE~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_DONE .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_DONE .power_up = "low";

cycloneive_lcell_comb \val_out~1 (
	.dataa(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datab(\fft_s2_cur.LPP_DONE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\val_out~1_combout ),
	.cout());
defparam \val_out~1 .lut_mask = 16'hEEEE;
defparam \val_out~1 .sum_lutc_input = "datac";

dffeas sop_out(
	.clk(clk),
	.d(\sop_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sop_out~q ),
	.prn(vcc));
defparam sop_out.is_wysiwyg = "true";
defparam sop_out.power_up = "low";

cycloneive_lcell_comb \master_source_sop~0 (
	.dataa(reset_n),
	.datab(\oe~q ),
	.datac(\sop_out~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\master_source_sop~0_combout ),
	.cout());
defparam \master_source_sop~0 .lut_mask = 16'hFEFE;
defparam \master_source_sop~0 .sum_lutc_input = "datac";

dffeas inv_i(
	.clk(clk),
	.d(\inv_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\inv_i~q ),
	.prn(vcc));
defparam inv_i.is_wysiwyg = "true";
defparam inv_i.power_up = "low";

cycloneive_lcell_comb \fft_dirn~0 (
	.dataa(\fft_dirn~q ),
	.datab(\inv_i~q ),
	.datac(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(\global_clock_enable~1_combout ),
	.cin(gnd),
	.combout(\fft_dirn~0_combout ),
	.cout());
defparam \fft_dirn~0 .lut_mask = 16'hEFFE;
defparam \fft_dirn~0 .sum_lutc_input = "datac";

dffeas exp_en(
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\exp_en~q ),
	.prn(vcc));
defparam exp_en.is_wysiwyg = "true";
defparam exp_en.power_up = "low";

cycloneive_lcell_comb \fft_s1_cur.NO_WRITE~5 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.DONE_WRITING~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s1_cur.NO_WRITE~5_combout ),
	.cout());
defparam \fft_s1_cur.NO_WRITE~5 .lut_mask = 16'hEEEE;
defparam \fft_s1_cur.NO_WRITE~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.DONE_WRITING~0 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.EARLY_DONE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s1_cur.DONE_WRITING~0_combout ),
	.cout());
defparam \fft_s1_cur.DONE_WRITING~0 .lut_mask = 16'hEEEE;
defparam \fft_s1_cur.DONE_WRITING~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.EARLY_DONE~0 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s1_cur.EARLY_DONE~0_combout ),
	.cout());
defparam \fft_s1_cur.EARLY_DONE~0 .lut_mask = 16'hEEEE;
defparam \fft_s1_cur.EARLY_DONE~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.FFT_PROCESS_A~0 (
	.dataa(reset_n),
	.datab(\fft_s1_cur.NO_WRITE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s1_cur.FFT_PROCESS_A~0_combout ),
	.cout());
defparam \fft_s1_cur.FFT_PROCESS_A~0 .lut_mask = 16'hEEEE;
defparam \fft_s1_cur.FFT_PROCESS_A~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \eop_out~0 (
	.dataa(\fft_s2_cur.START_LPP~q ),
	.datab(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datad(\bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ),
	.cin(gnd),
	.combout(\eop_out~0_combout ),
	.cout());
defparam \eop_out~0 .lut_mask = 16'hFF7F;
defparam \eop_out~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[23] (
	.clk(clk),
	.d(\data_rdy_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[23]~q ),
	.prn(vcc));
defparam \data_rdy_vec[23] .is_wysiwyg = "true";
defparam \data_rdy_vec[23] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~0 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~0_combout ),
	.cout());
defparam \data_rdy_vec~0 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.START_LPP~0 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\fft_s2_cur.START_LPP~0_combout ),
	.cout());
defparam \fft_s2_cur.START_LPP~0 .lut_mask = 16'hFEFE;
defparam \fft_s2_cur.START_LPP~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.WAIT_FOR_LPP_INPUT~0 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datac(\gen_radix_4_last_pass:lpp|gen_burst_val:delay_val|tdl_arr[4]~q ),
	.datad(\fft_s2_cur.START_LPP~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.WAIT_FOR_LPP_INPUT~0_combout ),
	.cout());
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~0 .lut_mask = 16'hFFBE;
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.WAIT_FOR_LPP_INPUT~1 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~0_combout ),
	.datab(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datac(\global_clock_enable~0_combout ),
	.datad(\auk_dsp_interface_controller_1|stall_reg~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.WAIT_FOR_LPP_INPUT~1_combout ),
	.cout());
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~1 .lut_mask = 16'hF737;
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.WAIT_FOR_LPP_INPUT~2 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.LPP_DONE~q ),
	.datac(\bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ),
	.datad(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.WAIT_FOR_LPP_INPUT~2_combout ),
	.cout());
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~2 .lut_mask = 16'hEFFF;
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.WAIT_FOR_LPP_INPUT~3 (
	.dataa(\fft_s2_cur.WAIT_FOR_LPP_INPUT~2_combout ),
	.datab(reset_n),
	.datac(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datad(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.WAIT_FOR_LPP_INPUT~3_combout ),
	.cout());
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~3 .lut_mask = 16'hFEFF;
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.LPP_OUTPUT_RDY~0 (
	.dataa(reset_n),
	.datab(\gen_radix_4_last_pass:lpp|gen_burst_val:delay_val|tdl_arr[4]~q ),
	.datac(\fft_s2_cur.START_LPP~q ),
	.datad(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.LPP_OUTPUT_RDY~0_combout ),
	.cout());
defparam \fft_s2_cur.LPP_OUTPUT_RDY~0 .lut_mask = 16'hFFFE;
defparam \fft_s2_cur.LPP_OUTPUT_RDY~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s2_cur.LPP_DONE~0 (
	.dataa(reset_n),
	.datab(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datac(gnd),
	.datad(\gen_radix_4_last_pass:lpp|gen_burst_val:delay_val|tdl_arr[4]~q ),
	.cin(gnd),
	.combout(\fft_s2_cur.LPP_DONE~0_combout ),
	.cout());
defparam \fft_s2_cur.LPP_DONE~0 .lut_mask = 16'hEEFF;
defparam \fft_s2_cur.LPP_DONE~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_out~0 (
	.dataa(\delay_sop|tdl_arr[6]~q ),
	.datab(\fft_s2_cur.START_LPP~q ),
	.datac(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sop_out~0_combout ),
	.cout());
defparam \sop_out~0 .lut_mask = 16'hFEFE;
defparam \sop_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_out~1 (
	.dataa(\sop_out~q ),
	.datab(\fft_s2_cur.START_LPP~q ),
	.datac(\fft_s2_cur.LPP_OUTPUT_RDY~q ),
	.datad(\fft_s2_cur.LPP_DONE~q ),
	.cin(gnd),
	.combout(\sop_out~1_combout ),
	.cout());
defparam \sop_out~1 .lut_mask = 16'hBFFF;
defparam \sop_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_out~2 (
	.dataa(\bfpdft|gen_disc:bfp_detect|sdetd.IDLE~q ),
	.datab(\sop_out~0_combout ),
	.datac(\sop_out~1_combout ),
	.datad(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.cin(gnd),
	.combout(\sop_out~2_combout ),
	.cout());
defparam \sop_out~2 .lut_mask = 16'hFEFF;
defparam \sop_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \inv_i~0 (
	.dataa(inverse_0),
	.datab(\inv_i~q ),
	.datac(gnd),
	.datad(sink_valid),
	.cin(gnd),
	.combout(\inv_i~0_combout ),
	.cout());
defparam \inv_i~0 .lut_mask = 16'hAACC;
defparam \inv_i~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[22] (
	.clk(clk),
	.d(\data_rdy_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[22]~q ),
	.prn(vcc));
defparam \data_rdy_vec[22] .is_wysiwyg = "true";
defparam \data_rdy_vec[22] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~1 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~1_combout ),
	.cout());
defparam \data_rdy_vec~1 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~1 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[21] (
	.clk(clk),
	.d(\data_rdy_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[21]~q ),
	.prn(vcc));
defparam \data_rdy_vec[21] .is_wysiwyg = "true";
defparam \data_rdy_vec[21] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~2 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~2_combout ),
	.cout());
defparam \data_rdy_vec~2 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~2 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[20] (
	.clk(clk),
	.d(\data_rdy_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[20]~q ),
	.prn(vcc));
defparam \data_rdy_vec[20] .is_wysiwyg = "true";
defparam \data_rdy_vec[20] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~3 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~3_combout ),
	.cout());
defparam \data_rdy_vec~3 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~3 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[19] (
	.clk(clk),
	.d(\data_rdy_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[19]~q ),
	.prn(vcc));
defparam \data_rdy_vec[19] .is_wysiwyg = "true";
defparam \data_rdy_vec[19] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~4 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~4_combout ),
	.cout());
defparam \data_rdy_vec~4 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~4 .sum_lutc_input = "datac";

dffeas \lpp_ram_data_out[3][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][12] .power_up = "low";

dffeas \lpp_ram_data_out[0][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][12] .power_up = "low";

dffeas \lpp_ram_data_out[1][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][12] .power_up = "low";

dffeas \lpp_ram_data_out[2][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][12] .power_up = "low";

dffeas \lpp_ram_data_out[3][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][2] .power_up = "low";

dffeas \lpp_ram_data_out[0][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][2] .power_up = "low";

dffeas \lpp_ram_data_out[1][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][2] .power_up = "low";

dffeas \lpp_ram_data_out[2][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][2] .power_up = "low";

dffeas \lpp_ram_data_out[3][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][11] .power_up = "low";

dffeas \lpp_ram_data_out[0][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][11] .power_up = "low";

dffeas \lpp_ram_data_out[1][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][11] .power_up = "low";

dffeas \lpp_ram_data_out[2][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][11] .power_up = "low";

dffeas \lpp_ram_data_out[3][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][1] .power_up = "low";

dffeas \lpp_ram_data_out[0][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][1] .power_up = "low";

dffeas \lpp_ram_data_out[1][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][1] .power_up = "low";

dffeas \lpp_ram_data_out[2][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][1] .power_up = "low";

dffeas \lpp_ram_data_out[3][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][10] .power_up = "low";

dffeas \lpp_ram_data_out[0][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][10] .power_up = "low";

dffeas \lpp_ram_data_out[1][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][10] .power_up = "low";

dffeas \lpp_ram_data_out[2][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][10] .power_up = "low";

dffeas \lpp_ram_data_out[3][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][0] .power_up = "low";

dffeas \lpp_ram_data_out[0][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][0] .power_up = "low";

dffeas \lpp_ram_data_out[1][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][0] .power_up = "low";

dffeas \lpp_ram_data_out[2][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][0] .power_up = "low";

dffeas \lpp_ram_data_out[3][19] (
	.clk(clk),
	.d(\lpp_ram_data_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][19]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][19] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][19] .power_up = "low";

dffeas \lpp_ram_data_out[0][19] (
	.clk(clk),
	.d(\lpp_ram_data_out~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][19]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][19] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][19] .power_up = "low";

dffeas \lpp_ram_data_out[1][19] (
	.clk(clk),
	.d(\lpp_ram_data_out~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][19]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][19] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][19] .power_up = "low";

dffeas \lpp_ram_data_out[2][19] (
	.clk(clk),
	.d(\lpp_ram_data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][19]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][19] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][19] .power_up = "low";

dffeas \lpp_ram_data_out[3][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][9] .power_up = "low";

dffeas \lpp_ram_data_out[0][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][9] .power_up = "low";

dffeas \lpp_ram_data_out[1][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][9] .power_up = "low";

dffeas \lpp_ram_data_out[2][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][9] .power_up = "low";

dffeas \lpp_ram_data_out[3][18] (
	.clk(clk),
	.d(\lpp_ram_data_out~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][18]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][18] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][18] .power_up = "low";

dffeas \lpp_ram_data_out[0][18] (
	.clk(clk),
	.d(\lpp_ram_data_out~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][18]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][18] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][18] .power_up = "low";

dffeas \lpp_ram_data_out[1][18] (
	.clk(clk),
	.d(\lpp_ram_data_out~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][18]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][18] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][18] .power_up = "low";

dffeas \lpp_ram_data_out[2][18] (
	.clk(clk),
	.d(\lpp_ram_data_out~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][18]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][18] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][18] .power_up = "low";

dffeas \lpp_ram_data_out[3][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][8] .power_up = "low";

dffeas \lpp_ram_data_out[0][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][8] .power_up = "low";

dffeas \lpp_ram_data_out[1][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][8] .power_up = "low";

dffeas \lpp_ram_data_out[2][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][8] .power_up = "low";

dffeas \lpp_ram_data_out[3][17] (
	.clk(clk),
	.d(\lpp_ram_data_out~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][17]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][17] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][17] .power_up = "low";

dffeas \lpp_ram_data_out[0][17] (
	.clk(clk),
	.d(\lpp_ram_data_out~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][17]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][17] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][17] .power_up = "low";

dffeas \lpp_ram_data_out[1][17] (
	.clk(clk),
	.d(\lpp_ram_data_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][17]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][17] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][17] .power_up = "low";

dffeas \lpp_ram_data_out[2][17] (
	.clk(clk),
	.d(\lpp_ram_data_out~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][17]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][17] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][17] .power_up = "low";

dffeas \lpp_ram_data_out[3][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][7] .power_up = "low";

dffeas \lpp_ram_data_out[0][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][7] .power_up = "low";

dffeas \lpp_ram_data_out[1][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][7] .power_up = "low";

dffeas \lpp_ram_data_out[2][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][7] .power_up = "low";

dffeas \lpp_ram_data_out[3][16] (
	.clk(clk),
	.d(\lpp_ram_data_out~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][16]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][16] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][16] .power_up = "low";

dffeas \lpp_ram_data_out[0][16] (
	.clk(clk),
	.d(\lpp_ram_data_out~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][16]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][16] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][16] .power_up = "low";

dffeas \lpp_ram_data_out[1][16] (
	.clk(clk),
	.d(\lpp_ram_data_out~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][16]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][16] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][16] .power_up = "low";

dffeas \lpp_ram_data_out[2][16] (
	.clk(clk),
	.d(\lpp_ram_data_out~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][16]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][16] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][16] .power_up = "low";

dffeas \lpp_ram_data_out[3][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][6] .power_up = "low";

dffeas \lpp_ram_data_out[0][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][6] .power_up = "low";

dffeas \lpp_ram_data_out[1][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][6] .power_up = "low";

dffeas \lpp_ram_data_out[2][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][6] .power_up = "low";

dffeas \lpp_ram_data_out[3][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][15] .power_up = "low";

dffeas \lpp_ram_data_out[0][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][15] .power_up = "low";

dffeas \lpp_ram_data_out[1][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][15] .power_up = "low";

dffeas \lpp_ram_data_out[2][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][15] .power_up = "low";

dffeas \lpp_ram_data_out[3][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][5] .power_up = "low";

dffeas \lpp_ram_data_out[0][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][5] .power_up = "low";

dffeas \lpp_ram_data_out[1][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][5] .power_up = "low";

dffeas \lpp_ram_data_out[2][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][5] .power_up = "low";

dffeas \lpp_ram_data_out[3][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][14] .power_up = "low";

dffeas \lpp_ram_data_out[0][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][14] .power_up = "low";

dffeas \lpp_ram_data_out[1][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][14] .power_up = "low";

dffeas \lpp_ram_data_out[2][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][14] .power_up = "low";

dffeas \lpp_ram_data_out[3][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][4] .power_up = "low";

dffeas \lpp_ram_data_out[0][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][4] .power_up = "low";

dffeas \lpp_ram_data_out[1][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][4] .power_up = "low";

dffeas \lpp_ram_data_out[2][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][4] .power_up = "low";

dffeas \lpp_ram_data_out[3][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][13] .power_up = "low";

dffeas \lpp_ram_data_out[0][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][13] .power_up = "low";

dffeas \lpp_ram_data_out[1][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][13] .power_up = "low";

dffeas \lpp_ram_data_out[2][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][13] .power_up = "low";

dffeas \lpp_ram_data_out[3][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[3][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][3] .power_up = "low";

dffeas \lpp_ram_data_out[0][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[0][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][3] .power_up = "low";

dffeas \lpp_ram_data_out[1][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[1][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][3] .power_up = "low";

dffeas \lpp_ram_data_out[2][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_ram_data_out[2][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][3] .power_up = "low";

dffeas \data_rdy_vec[18] (
	.clk(clk),
	.d(\data_rdy_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[18]~q ),
	.prn(vcc));
defparam \data_rdy_vec[18] .is_wysiwyg = "true";
defparam \data_rdy_vec[18] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~5 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~5_combout ),
	.cout());
defparam \data_rdy_vec~5 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~5 .sum_lutc_input = "datac";

dffeas \lpp_c_en_vec[6] (
	.clk(clk),
	.d(\lpp_c_en_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[6]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[6] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[6] .power_up = "low";

dffeas \lpp_c_en_vec[1] (
	.clk(clk),
	.d(\lpp_c_en_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[1]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[1] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[1] .power_up = "low";

cycloneive_lcell_comb \lpp_ram_data_out~0 (
	.dataa(reset_n),
	.datab(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datac(\lpp_c_en_vec[6]~q ),
	.datad(\lpp_c_en_vec[1]~q ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~0_combout ),
	.cout());
defparam \lpp_ram_data_out~0 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~1 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~1_combout ),
	.cout());
defparam \lpp_ram_data_out~1 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~2 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~2_combout ),
	.cout());
defparam \lpp_ram_data_out~2 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~3 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~3_combout ),
	.cout());
defparam \lpp_ram_data_out~3 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~4 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~4_combout ),
	.cout());
defparam \lpp_ram_data_out~4 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~5 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~5_combout ),
	.cout());
defparam \lpp_ram_data_out~5 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~6 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~6_combout ),
	.cout());
defparam \lpp_ram_data_out~6 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~7 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~7_combout ),
	.cout());
defparam \lpp_ram_data_out~7 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~8 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~8_combout ),
	.cout());
defparam \lpp_ram_data_out~8 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~9 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~9_combout ),
	.cout());
defparam \lpp_ram_data_out~9 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~10 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~10_combout ),
	.cout());
defparam \lpp_ram_data_out~10 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~11 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~11_combout ),
	.cout());
defparam \lpp_ram_data_out~11 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~12 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~12_combout ),
	.cout());
defparam \lpp_ram_data_out~12 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~13 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~13_combout ),
	.cout());
defparam \lpp_ram_data_out~13 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~14 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~14_combout ),
	.cout());
defparam \lpp_ram_data_out~14 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~15 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~15_combout ),
	.cout());
defparam \lpp_ram_data_out~15 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~16 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~16_combout ),
	.cout());
defparam \lpp_ram_data_out~16 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~17 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~17_combout ),
	.cout());
defparam \lpp_ram_data_out~17 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~18 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~18_combout ),
	.cout());
defparam \lpp_ram_data_out~18 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~19 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~19_combout ),
	.cout());
defparam \lpp_ram_data_out~19 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~20 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~20_combout ),
	.cout());
defparam \lpp_ram_data_out~20 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~21 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~21_combout ),
	.cout());
defparam \lpp_ram_data_out~21 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~22 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~22_combout ),
	.cout());
defparam \lpp_ram_data_out~22 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~23 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~23_combout ),
	.cout());
defparam \lpp_ram_data_out~23 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~24 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~24_combout ),
	.cout());
defparam \lpp_ram_data_out~24 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~25 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~25_combout ),
	.cout());
defparam \lpp_ram_data_out~25 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~26 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~26_combout ),
	.cout());
defparam \lpp_ram_data_out~26 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~27 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[19] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~27_combout ),
	.cout());
defparam \lpp_ram_data_out~27 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~28 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~28_combout ),
	.cout());
defparam \lpp_ram_data_out~28 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~29 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~29_combout ),
	.cout());
defparam \lpp_ram_data_out~29 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~30 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~30_combout ),
	.cout());
defparam \lpp_ram_data_out~30 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~31 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~31_combout ),
	.cout());
defparam \lpp_ram_data_out~31 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~32 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~32_combout ),
	.cout());
defparam \lpp_ram_data_out~32 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~33 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~33_combout ),
	.cout());
defparam \lpp_ram_data_out~33 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~34 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~34_combout ),
	.cout());
defparam \lpp_ram_data_out~34 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~35 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[18] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~35_combout ),
	.cout());
defparam \lpp_ram_data_out~35 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~36 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~36_combout ),
	.cout());
defparam \lpp_ram_data_out~36 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~37 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~37_combout ),
	.cout());
defparam \lpp_ram_data_out~37 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~38 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~38_combout ),
	.cout());
defparam \lpp_ram_data_out~38 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~39 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~39_combout ),
	.cout());
defparam \lpp_ram_data_out~39 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~40 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~40_combout ),
	.cout());
defparam \lpp_ram_data_out~40 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~41 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~41_combout ),
	.cout());
defparam \lpp_ram_data_out~41 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~42 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~42_combout ),
	.cout());
defparam \lpp_ram_data_out~42 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~43 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[17] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~43_combout ),
	.cout());
defparam \lpp_ram_data_out~43 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~44 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~44_combout ),
	.cout());
defparam \lpp_ram_data_out~44 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~45 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~45_combout ),
	.cout());
defparam \lpp_ram_data_out~45 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~46 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~46_combout ),
	.cout());
defparam \lpp_ram_data_out~46 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~47 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~47_combout ),
	.cout());
defparam \lpp_ram_data_out~47 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~48 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~48_combout ),
	.cout());
defparam \lpp_ram_data_out~48 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~49 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~49_combout ),
	.cout());
defparam \lpp_ram_data_out~49 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~50 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~50_combout ),
	.cout());
defparam \lpp_ram_data_out~50 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~51 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[16] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~51_combout ),
	.cout());
defparam \lpp_ram_data_out~51 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~52 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~52_combout ),
	.cout());
defparam \lpp_ram_data_out~52 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~53 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~53_combout ),
	.cout());
defparam \lpp_ram_data_out~53 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~54 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~54_combout ),
	.cout());
defparam \lpp_ram_data_out~54 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~55 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~55_combout ),
	.cout());
defparam \lpp_ram_data_out~55 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~56 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~56_combout ),
	.cout());
defparam \lpp_ram_data_out~56 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~57 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~57_combout ),
	.cout());
defparam \lpp_ram_data_out~57 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~58 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~58_combout ),
	.cout());
defparam \lpp_ram_data_out~58 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~59 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~59_combout ),
	.cout());
defparam \lpp_ram_data_out~59 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~60 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~60_combout ),
	.cout());
defparam \lpp_ram_data_out~60 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~61 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~61_combout ),
	.cout());
defparam \lpp_ram_data_out~61 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~62 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~62_combout ),
	.cout());
defparam \lpp_ram_data_out~62 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~63 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~63_combout ),
	.cout());
defparam \lpp_ram_data_out~63 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~64 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~64_combout ),
	.cout());
defparam \lpp_ram_data_out~64 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~65 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~65_combout ),
	.cout());
defparam \lpp_ram_data_out~65 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~66 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~66_combout ),
	.cout());
defparam \lpp_ram_data_out~66 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~67 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~67_combout ),
	.cout());
defparam \lpp_ram_data_out~67 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~68 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~68_combout ),
	.cout());
defparam \lpp_ram_data_out~68 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~69 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~69_combout ),
	.cout());
defparam \lpp_ram_data_out~69 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~70 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~70_combout ),
	.cout());
defparam \lpp_ram_data_out~70 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~71 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~71_combout ),
	.cout());
defparam \lpp_ram_data_out~71 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~72 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~72_combout ),
	.cout());
defparam \lpp_ram_data_out~72 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~73 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~73_combout ),
	.cout());
defparam \lpp_ram_data_out~73 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~74 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~74_combout ),
	.cout());
defparam \lpp_ram_data_out~74 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~75 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~75_combout ),
	.cout());
defparam \lpp_ram_data_out~75 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~76 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~76_combout ),
	.cout());
defparam \lpp_ram_data_out~76 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~77 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~77_combout ),
	.cout());
defparam \lpp_ram_data_out~77 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~78 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~78_combout ),
	.cout());
defparam \lpp_ram_data_out~78 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_ram_data_out~79 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[6]~q ),
	.datac(\lpp_c_en_vec[1]~q ),
	.datad(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.cin(gnd),
	.combout(\lpp_ram_data_out~79_combout ),
	.cout());
defparam \lpp_ram_data_out~79 .lut_mask = 16'hFFFE;
defparam \lpp_ram_data_out~79 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[17] (
	.clk(clk),
	.d(\data_rdy_vec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[17]~q ),
	.prn(vcc));
defparam \data_rdy_vec[17] .is_wysiwyg = "true";
defparam \data_rdy_vec[17] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~6 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~6_combout ),
	.cout());
defparam \data_rdy_vec~6 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~6 .sum_lutc_input = "datac";

dffeas \wren_a[3] (
	.clk(clk),
	.d(\wren_a~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wren_a[3]~q ),
	.prn(vcc));
defparam \wren_a[3] .is_wysiwyg = "true";
defparam \wren_a[3] .power_up = "low";

dffeas \lpp_c_en_vec[5] (
	.clk(clk),
	.d(\lpp_c_en_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[5]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[5] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[5] .power_up = "low";

cycloneive_lcell_comb \lpp_c_en_vec~0 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~0_combout ),
	.cout());
defparam \lpp_c_en_vec~0 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_c_en_vec~1 (
	.dataa(reset_n),
	.datab(\gen_radix_4_last_pass:gen_lpp_addr|en_d~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~1_combout ),
	.cout());
defparam \lpp_c_en_vec~1 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~1 .sum_lutc_input = "datac";

dffeas \wren_a[0] (
	.clk(clk),
	.d(\wren_a~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wren_a[0]~q ),
	.prn(vcc));
defparam \wren_a[0] .is_wysiwyg = "true";
defparam \wren_a[0] .power_up = "low";

dffeas \wren_a[1] (
	.clk(clk),
	.d(\wren_a~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wren_a[1]~q ),
	.prn(vcc));
defparam \wren_a[1] .is_wysiwyg = "true";
defparam \wren_a[1] .power_up = "low";

dffeas \wren_a[2] (
	.clk(clk),
	.d(\wren_a~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wren_a[2]~q ),
	.prn(vcc));
defparam \wren_a[2] .is_wysiwyg = "true";
defparam \wren_a[2] .power_up = "low";

dffeas \data_rdy_vec[16] (
	.clk(clk),
	.d(\data_rdy_vec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[16]~q ),
	.prn(vcc));
defparam \data_rdy_vec[16] .is_wysiwyg = "true";
defparam \data_rdy_vec[16] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~7 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~7_combout ),
	.cout());
defparam \data_rdy_vec~7 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~7 .sum_lutc_input = "datac";

dffeas \wc_vec[3] (
	.clk(clk),
	.d(\wc_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wc_vec[3]~q ),
	.prn(vcc));
defparam \wc_vec[3] .is_wysiwyg = "true";
defparam \wc_vec[3] .power_up = "low";

cycloneive_lcell_comb \wren_a~2 (
	.dataa(\fft_s1_cur.WAIT_FOR_INPUT~0_combout ),
	.datab(\wc_vec[3]~q ),
	.datac(\writer|data_rdy_int~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\wren_a~2_combout ),
	.cout());
defparam \wren_a~2 .lut_mask = 16'hFEFE;
defparam \wren_a~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_s1_cur.WAIT_FOR_INPUT~4 (
	.dataa(gnd),
	.datab(\fft_s1_cur.WRITE_INPUT~q ),
	.datac(\fft_s1_cur.DONE_WRITING~q ),
	.datad(\fft_s1_cur.EARLY_DONE~q ),
	.cin(gnd),
	.combout(\fft_s1_cur.WAIT_FOR_INPUT~4_combout ),
	.cout());
defparam \fft_s1_cur.WAIT_FOR_INPUT~4 .lut_mask = 16'h3FFF;
defparam \fft_s1_cur.WAIT_FOR_INPUT~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wren_a~3 (
	.dataa(\fft_s1_cur.IDLE~q ),
	.datab(\wren_a~2_combout ),
	.datac(\writer|wren[3]~q ),
	.datad(\fft_s1_cur.WAIT_FOR_INPUT~4_combout ),
	.cin(gnd),
	.combout(\wren_a~3_combout ),
	.cout());
defparam \wren_a~3 .lut_mask = 16'hFEFF;
defparam \wren_a~3 .sum_lutc_input = "datac";

dffeas sel_ram_in(
	.clk(clk),
	.d(\sel_ram_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sel_ram_in~q ),
	.prn(vcc));
defparam sel_ram_in.is_wysiwyg = "true";
defparam sel_ram_in.power_up = "low";

dffeas \data_rdy_vec[2] (
	.clk(clk),
	.d(\data_rdy_vec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[2]~q ),
	.prn(vcc));
defparam \data_rdy_vec[2] .is_wysiwyg = "true";
defparam \data_rdy_vec[2] .power_up = "low";

dffeas \data_rdy_vec[0] (
	.clk(clk),
	.d(\data_rdy_vec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[0]~q ),
	.prn(vcc));
defparam \data_rdy_vec[0] .is_wysiwyg = "true";
defparam \data_rdy_vec[0] .power_up = "low";

dffeas \lpp_c_en_vec[4] (
	.clk(clk),
	.d(\lpp_c_en_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[4]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[4] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[4] .power_up = "low";

cycloneive_lcell_comb \lpp_c_en_vec~2 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~2_combout ),
	.cout());
defparam \lpp_c_en_vec~2 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wren_a~4 (
	.dataa(\fft_s1_cur.IDLE~q ),
	.datab(\wren_a~2_combout ),
	.datac(\writer|wren[0]~q ),
	.datad(\fft_s1_cur.WAIT_FOR_INPUT~4_combout ),
	.cin(gnd),
	.combout(\wren_a~4_combout ),
	.cout());
defparam \wren_a~4 .lut_mask = 16'hFEFF;
defparam \wren_a~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wren_a~5 (
	.dataa(\fft_s1_cur.IDLE~q ),
	.datab(\wren_a~2_combout ),
	.datac(\writer|wren[1]~q ),
	.datad(\fft_s1_cur.WAIT_FOR_INPUT~4_combout ),
	.cin(gnd),
	.combout(\wren_a~5_combout ),
	.cout());
defparam \wren_a~5 .lut_mask = 16'hFEFF;
defparam \wren_a~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wren_a~6 (
	.dataa(\fft_s1_cur.IDLE~q ),
	.datab(\wren_a~2_combout ),
	.datac(\writer|wren[2]~q ),
	.datad(\fft_s1_cur.WAIT_FOR_INPUT~4_combout ),
	.cin(gnd),
	.combout(\wren_a~6_combout ),
	.cout());
defparam \wren_a~6 .lut_mask = 16'hFEFF;
defparam \wren_a~6 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[15] (
	.clk(clk),
	.d(\data_rdy_vec~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[15]~q ),
	.prn(vcc));
defparam \data_rdy_vec[15] .is_wysiwyg = "true";
defparam \data_rdy_vec[15] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~8 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~8_combout ),
	.cout());
defparam \data_rdy_vec~8 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~8 .sum_lutc_input = "datac";

dffeas \wc_vec[2] (
	.clk(clk),
	.d(\wc_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wc_vec[2]~q ),
	.prn(vcc));
defparam \wc_vec[2] .is_wysiwyg = "true";
defparam \wc_vec[2] .power_up = "low";

cycloneive_lcell_comb \wc_vec~0 (
	.dataa(reset_n),
	.datab(\wc_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~0_combout ),
	.cout());
defparam \wc_vec~0 .lut_mask = 16'hEEEE;
defparam \wc_vec~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sel_ram_in~0 (
	.dataa(\fft_s1_cur.WRITE_INPUT~q ),
	.datab(\fft_s1_cur.DONE_WRITING~q ),
	.datac(\fft_s1_cur.EARLY_DONE~q ),
	.datad(\fft_s1_cur.IDLE~q ),
	.cin(gnd),
	.combout(\sel_ram_in~0_combout ),
	.cout());
defparam \sel_ram_in~0 .lut_mask = 16'hFF7F;
defparam \sel_ram_in~0 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[1] (
	.clk(clk),
	.d(\data_rdy_vec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[1]~q ),
	.prn(vcc));
defparam \data_rdy_vec[1] .is_wysiwyg = "true";
defparam \data_rdy_vec[1] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~9 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~9_combout ),
	.cout());
defparam \data_rdy_vec~9 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~10 (
	.dataa(reset_n),
	.datab(\writer|data_rdy_int~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~10_combout ),
	.cout());
defparam \data_rdy_vec~10 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~10 .sum_lutc_input = "datac";

dffeas \lpp_c_en_vec[3] (
	.clk(clk),
	.d(\lpp_c_en_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[3]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[3] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[3] .power_up = "low";

cycloneive_lcell_comb \lpp_c_en_vec~3 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~3_combout ),
	.cout());
defparam \lpp_c_en_vec~3 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~3 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[14] (
	.clk(clk),
	.d(\data_rdy_vec~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[14]~q ),
	.prn(vcc));
defparam \data_rdy_vec[14] .is_wysiwyg = "true";
defparam \data_rdy_vec[14] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~11 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~11_combout ),
	.cout());
defparam \data_rdy_vec~11 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~11 .sum_lutc_input = "datac";

dffeas \p_cd_en[2] (
	.clk(clk),
	.d(\reg_we_window~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_cd_en[2]~q ),
	.prn(vcc));
defparam \p_cd_en[2] .is_wysiwyg = "true";
defparam \p_cd_en[2] .power_up = "low";

dffeas \wc_vec[1] (
	.clk(clk),
	.d(\wc_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\wc_vec[1]~q ),
	.prn(vcc));
defparam \wc_vec[1] .is_wysiwyg = "true";
defparam \wc_vec[1] .power_up = "low";

cycloneive_lcell_comb \wc_vec~1 (
	.dataa(reset_n),
	.datab(\wc_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~1_combout ),
	.cout());
defparam \wc_vec~1 .lut_mask = 16'hEEEE;
defparam \wc_vec~1 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[2] (
	.clk(clk),
	.d(\data_imag_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[2]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[2] .is_wysiwyg = "true";
defparam \data_imag_in_reg[2] .power_up = "low";

dffeas \data_real_in_reg[2] (
	.clk(clk),
	.d(\data_real_in_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[2]~q ),
	.prn(vcc));
defparam \data_real_in_reg[2] .is_wysiwyg = "true";
defparam \data_real_in_reg[2] .power_up = "low";

cycloneive_lcell_comb \core_real_in~0 (
	.dataa(\data_imag_in_reg[2]~q ),
	.datab(\data_real_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~0_combout ),
	.cout());
defparam \core_real_in~0 .lut_mask = 16'hAACC;
defparam \core_real_in~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~12 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~12_combout ),
	.cout());
defparam \data_rdy_vec~12 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~12 .sum_lutc_input = "datac";

dffeas \lpp_c_en_vec[2] (
	.clk(clk),
	.d(\lpp_c_en_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\lpp_c_en_vec[2]~q ),
	.prn(vcc));
defparam \lpp_c_en_vec[2] .is_wysiwyg = "true";
defparam \lpp_c_en_vec[2] .power_up = "low";

cycloneive_lcell_comb \lpp_c_en_vec~4 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~4_combout ),
	.cout());
defparam \lpp_c_en_vec~4 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~0 (
	.dataa(\data_real_in_reg[2]~q ),
	.datab(\data_imag_in_reg[2]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~0_combout ),
	.cout());
defparam \core_imag_in~0 .lut_mask = 16'hAACC;
defparam \core_imag_in~0 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[1] (
	.clk(clk),
	.d(\data_imag_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[1]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[1] .is_wysiwyg = "true";
defparam \data_imag_in_reg[1] .power_up = "low";

dffeas \data_real_in_reg[1] (
	.clk(clk),
	.d(\data_real_in_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[1]~q ),
	.prn(vcc));
defparam \data_real_in_reg[1] .is_wysiwyg = "true";
defparam \data_real_in_reg[1] .power_up = "low";

cycloneive_lcell_comb \core_real_in~1 (
	.dataa(\data_imag_in_reg[1]~q ),
	.datab(\data_real_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~1_combout ),
	.cout());
defparam \core_real_in~1 .lut_mask = 16'hAACC;
defparam \core_real_in~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~1 (
	.dataa(\data_real_in_reg[1]~q ),
	.datab(\data_imag_in_reg[1]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~1_combout ),
	.cout());
defparam \core_imag_in~1 .lut_mask = 16'hAACC;
defparam \core_imag_in~1 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[0] (
	.clk(clk),
	.d(\data_imag_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[0]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[0] .is_wysiwyg = "true";
defparam \data_imag_in_reg[0] .power_up = "low";

dffeas \data_real_in_reg[0] (
	.clk(clk),
	.d(\data_real_in_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[0]~q ),
	.prn(vcc));
defparam \data_real_in_reg[0] .is_wysiwyg = "true";
defparam \data_real_in_reg[0] .power_up = "low";

cycloneive_lcell_comb \core_real_in~2 (
	.dataa(\data_imag_in_reg[0]~q ),
	.datab(\data_real_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~2_combout ),
	.cout());
defparam \core_real_in~2 .lut_mask = 16'hAACC;
defparam \core_real_in~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~2 (
	.dataa(\data_real_in_reg[0]~q ),
	.datab(\data_imag_in_reg[0]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~2_combout ),
	.cout());
defparam \core_imag_in~2 .lut_mask = 16'hAACC;
defparam \core_imag_in~2 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[9] (
	.clk(clk),
	.d(\data_imag_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[9]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[9] .is_wysiwyg = "true";
defparam \data_imag_in_reg[9] .power_up = "low";

dffeas \data_real_in_reg[9] (
	.clk(clk),
	.d(\data_real_in_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[9]~q ),
	.prn(vcc));
defparam \data_real_in_reg[9] .is_wysiwyg = "true";
defparam \data_real_in_reg[9] .power_up = "low";

cycloneive_lcell_comb \core_real_in~3 (
	.dataa(\data_imag_in_reg[9]~q ),
	.datab(\data_real_in_reg[9]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~3_combout ),
	.cout());
defparam \core_real_in~3 .lut_mask = 16'hAACC;
defparam \core_real_in~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~3 (
	.dataa(\data_real_in_reg[9]~q ),
	.datab(\data_imag_in_reg[9]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~3_combout ),
	.cout());
defparam \core_imag_in~3 .lut_mask = 16'hAACC;
defparam \core_imag_in~3 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[8] (
	.clk(clk),
	.d(\data_imag_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[8]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[8] .is_wysiwyg = "true";
defparam \data_imag_in_reg[8] .power_up = "low";

dffeas \data_real_in_reg[8] (
	.clk(clk),
	.d(\data_real_in_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[8]~q ),
	.prn(vcc));
defparam \data_real_in_reg[8] .is_wysiwyg = "true";
defparam \data_real_in_reg[8] .power_up = "low";

cycloneive_lcell_comb \core_real_in~4 (
	.dataa(\data_imag_in_reg[8]~q ),
	.datab(\data_real_in_reg[8]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~4_combout ),
	.cout());
defparam \core_real_in~4 .lut_mask = 16'hAACC;
defparam \core_real_in~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~4 (
	.dataa(\data_real_in_reg[8]~q ),
	.datab(\data_imag_in_reg[8]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~4_combout ),
	.cout());
defparam \core_imag_in~4 .lut_mask = 16'hAACC;
defparam \core_imag_in~4 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[7] (
	.clk(clk),
	.d(\data_imag_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[7]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[7] .is_wysiwyg = "true";
defparam \data_imag_in_reg[7] .power_up = "low";

dffeas \data_real_in_reg[7] (
	.clk(clk),
	.d(\data_real_in_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[7]~q ),
	.prn(vcc));
defparam \data_real_in_reg[7] .is_wysiwyg = "true";
defparam \data_real_in_reg[7] .power_up = "low";

cycloneive_lcell_comb \core_real_in~5 (
	.dataa(\data_imag_in_reg[7]~q ),
	.datab(\data_real_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~5_combout ),
	.cout());
defparam \core_real_in~5 .lut_mask = 16'hAACC;
defparam \core_real_in~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~5 (
	.dataa(\data_real_in_reg[7]~q ),
	.datab(\data_imag_in_reg[7]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~5_combout ),
	.cout());
defparam \core_imag_in~5 .lut_mask = 16'hAACC;
defparam \core_imag_in~5 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[6] (
	.clk(clk),
	.d(\data_imag_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[6]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[6] .is_wysiwyg = "true";
defparam \data_imag_in_reg[6] .power_up = "low";

dffeas \data_real_in_reg[6] (
	.clk(clk),
	.d(\data_real_in_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[6]~q ),
	.prn(vcc));
defparam \data_real_in_reg[6] .is_wysiwyg = "true";
defparam \data_real_in_reg[6] .power_up = "low";

cycloneive_lcell_comb \core_real_in~6 (
	.dataa(\data_imag_in_reg[6]~q ),
	.datab(\data_real_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~6_combout ),
	.cout());
defparam \core_real_in~6 .lut_mask = 16'hAACC;
defparam \core_real_in~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~6 (
	.dataa(\data_real_in_reg[6]~q ),
	.datab(\data_imag_in_reg[6]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~6_combout ),
	.cout());
defparam \core_imag_in~6 .lut_mask = 16'hAACC;
defparam \core_imag_in~6 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[5] (
	.clk(clk),
	.d(\data_imag_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[5]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[5] .is_wysiwyg = "true";
defparam \data_imag_in_reg[5] .power_up = "low";

dffeas \data_real_in_reg[5] (
	.clk(clk),
	.d(\data_real_in_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[5]~q ),
	.prn(vcc));
defparam \data_real_in_reg[5] .is_wysiwyg = "true";
defparam \data_real_in_reg[5] .power_up = "low";

cycloneive_lcell_comb \core_real_in~7 (
	.dataa(\data_imag_in_reg[5]~q ),
	.datab(\data_real_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~7_combout ),
	.cout());
defparam \core_real_in~7 .lut_mask = 16'hAACC;
defparam \core_real_in~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~7 (
	.dataa(\data_real_in_reg[5]~q ),
	.datab(\data_imag_in_reg[5]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~7_combout ),
	.cout());
defparam \core_imag_in~7 .lut_mask = 16'hAACC;
defparam \core_imag_in~7 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[4] (
	.clk(clk),
	.d(\data_imag_in_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[4]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[4] .is_wysiwyg = "true";
defparam \data_imag_in_reg[4] .power_up = "low";

dffeas \data_real_in_reg[4] (
	.clk(clk),
	.d(\data_real_in_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[4]~q ),
	.prn(vcc));
defparam \data_real_in_reg[4] .is_wysiwyg = "true";
defparam \data_real_in_reg[4] .power_up = "low";

cycloneive_lcell_comb \core_real_in~8 (
	.dataa(\data_imag_in_reg[4]~q ),
	.datab(\data_real_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~8_combout ),
	.cout());
defparam \core_real_in~8 .lut_mask = 16'hAACC;
defparam \core_real_in~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~8 (
	.dataa(\data_real_in_reg[4]~q ),
	.datab(\data_imag_in_reg[4]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~8_combout ),
	.cout());
defparam \core_imag_in~8 .lut_mask = 16'hAACC;
defparam \core_imag_in~8 .sum_lutc_input = "datac";

dffeas \data_imag_in_reg[3] (
	.clk(clk),
	.d(\data_imag_in_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_imag_in_reg[3]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[3] .is_wysiwyg = "true";
defparam \data_imag_in_reg[3] .power_up = "low";

dffeas \data_real_in_reg[3] (
	.clk(clk),
	.d(\data_real_in_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_real_in_reg[3]~q ),
	.prn(vcc));
defparam \data_real_in_reg[3] .is_wysiwyg = "true";
defparam \data_real_in_reg[3] .power_up = "low";

cycloneive_lcell_comb \core_real_in~9 (
	.dataa(\data_imag_in_reg[3]~q ),
	.datab(\data_real_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_real_in~9_combout ),
	.cout());
defparam \core_real_in~9 .lut_mask = 16'hAACC;
defparam \core_real_in~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \core_imag_in~9 (
	.dataa(\data_real_in_reg[3]~q ),
	.datab(\data_imag_in_reg[3]~q ),
	.datac(gnd),
	.datad(\fft_dirn~q ),
	.cin(gnd),
	.combout(\core_imag_in~9_combout ),
	.cout());
defparam \core_imag_in~9 .lut_mask = 16'hAACC;
defparam \core_imag_in~9 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[13] (
	.clk(clk),
	.d(\data_rdy_vec~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[13]~q ),
	.prn(vcc));
defparam \data_rdy_vec[13] .is_wysiwyg = "true";
defparam \data_rdy_vec[13] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~13 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~13_combout ),
	.cout());
defparam \data_rdy_vec~13 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~13 .sum_lutc_input = "datac";

dffeas \p_tdl[13][2] (
	.clk(clk),
	.d(\p_tdl~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[13][2]~q ),
	.prn(vcc));
defparam \p_tdl[13][2] .is_wysiwyg = "true";
defparam \p_tdl[13][2] .power_up = "low";

dffeas \p_tdl[13][0] (
	.clk(clk),
	.d(\p_tdl~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[13][0]~q ),
	.prn(vcc));
defparam \p_tdl[13][0] .is_wysiwyg = "true";
defparam \p_tdl[13][0] .power_up = "low";

dffeas \p_tdl[13][1] (
	.clk(clk),
	.d(\p_tdl~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[13][1]~q ),
	.prn(vcc));
defparam \p_tdl[13][1] .is_wysiwyg = "true";
defparam \p_tdl[13][1] .power_up = "low";

dffeas \p_tdl[11][0] (
	.clk(clk),
	.d(\p_tdl~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[11][0]~q ),
	.prn(vcc));
defparam \p_tdl[11][0] .is_wysiwyg = "true";
defparam \p_tdl[11][0] .power_up = "low";

cycloneive_lcell_comb \reg_we_window~0 (
	.dataa(\p_tdl[13][2]~q ),
	.datab(\p_tdl[13][0]~q ),
	.datac(\p_tdl[13][1]~q ),
	.datad(\p_tdl[11][0]~q ),
	.cin(gnd),
	.combout(\reg_we_window~0_combout ),
	.cout());
defparam \reg_we_window~0 .lut_mask = 16'hBFFF;
defparam \reg_we_window~0 .sum_lutc_input = "datac";

dffeas \p_tdl[11][2] (
	.clk(clk),
	.d(\p_tdl~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[11][2]~q ),
	.prn(vcc));
defparam \p_tdl[11][2] .is_wysiwyg = "true";
defparam \p_tdl[11][2] .power_up = "low";

dffeas \p_tdl[11][1] (
	.clk(clk),
	.d(\p_tdl~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[11][1]~q ),
	.prn(vcc));
defparam \p_tdl[11][1] .is_wysiwyg = "true";
defparam \p_tdl[11][1] .power_up = "low";

cycloneive_lcell_comb \reg_we_window~1 (
	.dataa(\reg_we_window~0_combout ),
	.datab(\p_tdl[11][2]~q ),
	.datac(gnd),
	.datad(\p_tdl[11][1]~q ),
	.cin(gnd),
	.combout(\reg_we_window~1_combout ),
	.cout());
defparam \reg_we_window~1 .lut_mask = 16'hEEFF;
defparam \reg_we_window~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wc_vec~2 (
	.dataa(reset_n),
	.datab(\sel_we|wc_i_d~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_vec~2_combout ),
	.cout());
defparam \wc_vec~2 .lut_mask = 16'hEEEE;
defparam \wc_vec~2 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[4] (
	.clk(clk),
	.d(\data_rdy_vec~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[4]~q ),
	.prn(vcc));
defparam \data_rdy_vec[4] .is_wysiwyg = "true";
defparam \data_rdy_vec[4] .power_up = "low";

cycloneive_lcell_comb \data_imag_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~0_combout ),
	.cout());
defparam \data_imag_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~0 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~0_combout ),
	.cout());
defparam \data_real_in_reg~0 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \lpp_c_en_vec~5 (
	.dataa(reset_n),
	.datab(\lpp_c_en_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\lpp_c_en_vec~5_combout ),
	.cout());
defparam \lpp_c_en_vec~5 .lut_mask = 16'hEEEE;
defparam \lpp_c_en_vec~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~1_combout ),
	.cout());
defparam \data_imag_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~1 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~1_combout ),
	.cout());
defparam \data_real_in_reg~1 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~2_combout ),
	.cout());
defparam \data_imag_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~2 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~2_combout ),
	.cout());
defparam \data_real_in_reg~2 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~3_combout ),
	.cout());
defparam \data_imag_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~3 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~3_combout ),
	.cout());
defparam \data_real_in_reg~3 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~4_combout ),
	.cout());
defparam \data_imag_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~4 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~4_combout ),
	.cout());
defparam \data_real_in_reg~4 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~5_combout ),
	.cout());
defparam \data_imag_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~5 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~5_combout ),
	.cout());
defparam \data_real_in_reg~5 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~6_combout ),
	.cout());
defparam \data_imag_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~6 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~6_combout ),
	.cout());
defparam \data_real_in_reg~6 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~7_combout ),
	.cout());
defparam \data_imag_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~7 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~7_combout ),
	.cout());
defparam \data_real_in_reg~7 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~8 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~8_combout ),
	.cout());
defparam \data_imag_in_reg~8 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~8 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~8_combout ),
	.cout());
defparam \data_real_in_reg~8 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_imag_in_reg~9 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_imag_in_reg~9_combout ),
	.cout());
defparam \data_imag_in_reg~9 .lut_mask = 16'hEEEE;
defparam \data_imag_in_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_in_reg~9 (
	.dataa(reset_n),
	.datab(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_in_reg~9_combout ),
	.cout());
defparam \data_real_in_reg~9 .lut_mask = 16'hEEEE;
defparam \data_real_in_reg~9 .sum_lutc_input = "datac";

dffeas \twiddle_data[0][1][0] (
	.clk(clk),
	.d(\twiddle_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][0] .power_up = "low";

dffeas \twiddle_data[0][1][1] (
	.clk(clk),
	.d(\twiddle_data~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][1] .power_up = "low";

dffeas \twiddle_data[0][1][2] (
	.clk(clk),
	.d(\twiddle_data~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][2] .power_up = "low";

dffeas \twiddle_data[0][1][3] (
	.clk(clk),
	.d(\twiddle_data~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][3] .power_up = "low";

dffeas \twiddle_data[0][1][4] (
	.clk(clk),
	.d(\twiddle_data~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][4] .power_up = "low";

dffeas \twiddle_data[0][1][5] (
	.clk(clk),
	.d(\twiddle_data~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][5] .power_up = "low";

dffeas \twiddle_data[0][1][6] (
	.clk(clk),
	.d(\twiddle_data~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][6] .power_up = "low";

dffeas \twiddle_data[0][1][7] (
	.clk(clk),
	.d(\twiddle_data~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][7] .power_up = "low";

dffeas \twiddle_data[0][1][8] (
	.clk(clk),
	.d(\twiddle_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][8]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][8] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][8] .power_up = "low";

dffeas \twiddle_data[0][1][9] (
	.clk(clk),
	.d(\twiddle_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][1][9]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][9] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][9] .power_up = "low";

dffeas \twiddle_data[0][0][0] (
	.clk(clk),
	.d(\twiddle_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][0] .power_up = "low";

dffeas \twiddle_data[0][0][1] (
	.clk(clk),
	.d(\twiddle_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][1] .power_up = "low";

dffeas \twiddle_data[0][0][2] (
	.clk(clk),
	.d(\twiddle_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][2] .power_up = "low";

dffeas \twiddle_data[0][0][3] (
	.clk(clk),
	.d(\twiddle_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][3] .power_up = "low";

dffeas \twiddle_data[0][0][4] (
	.clk(clk),
	.d(\twiddle_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][4] .power_up = "low";

dffeas \twiddle_data[0][0][5] (
	.clk(clk),
	.d(\twiddle_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][5] .power_up = "low";

dffeas \twiddle_data[0][0][6] (
	.clk(clk),
	.d(\twiddle_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][6] .power_up = "low";

dffeas \twiddle_data[0][0][7] (
	.clk(clk),
	.d(\twiddle_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][7] .power_up = "low";

dffeas \twiddle_data[0][0][8] (
	.clk(clk),
	.d(\twiddle_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][8]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][8] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][8] .power_up = "low";

dffeas \twiddle_data[0][0][9] (
	.clk(clk),
	.d(\twiddle_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[0][0][9]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][9] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][9] .power_up = "low";

dffeas \twiddle_data[1][1][0] (
	.clk(clk),
	.d(\twiddle_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][0] .power_up = "low";

dffeas \twiddle_data[1][1][1] (
	.clk(clk),
	.d(\twiddle_data~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][1] .power_up = "low";

dffeas \twiddle_data[1][1][2] (
	.clk(clk),
	.d(\twiddle_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][2] .power_up = "low";

dffeas \twiddle_data[1][1][3] (
	.clk(clk),
	.d(\twiddle_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][3] .power_up = "low";

dffeas \twiddle_data[1][1][4] (
	.clk(clk),
	.d(\twiddle_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][4] .power_up = "low";

dffeas \twiddle_data[1][1][5] (
	.clk(clk),
	.d(\twiddle_data~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][5] .power_up = "low";

dffeas \twiddle_data[1][1][6] (
	.clk(clk),
	.d(\twiddle_data~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][6] .power_up = "low";

dffeas \twiddle_data[1][1][7] (
	.clk(clk),
	.d(\twiddle_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][7] .power_up = "low";

dffeas \twiddle_data[1][1][8] (
	.clk(clk),
	.d(\twiddle_data~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][8]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][8] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][8] .power_up = "low";

dffeas \twiddle_data[1][1][9] (
	.clk(clk),
	.d(\twiddle_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][1][9]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][9] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][9] .power_up = "low";

dffeas \twiddle_data[1][0][0] (
	.clk(clk),
	.d(\twiddle_data~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][0] .power_up = "low";

dffeas \twiddle_data[1][0][1] (
	.clk(clk),
	.d(\twiddle_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][1] .power_up = "low";

dffeas \twiddle_data[1][0][2] (
	.clk(clk),
	.d(\twiddle_data~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][2] .power_up = "low";

dffeas \twiddle_data[1][0][3] (
	.clk(clk),
	.d(\twiddle_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][3] .power_up = "low";

dffeas \twiddle_data[1][0][4] (
	.clk(clk),
	.d(\twiddle_data~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][4] .power_up = "low";

dffeas \twiddle_data[1][0][5] (
	.clk(clk),
	.d(\twiddle_data~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][5] .power_up = "low";

dffeas \twiddle_data[1][0][6] (
	.clk(clk),
	.d(\twiddle_data~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][6] .power_up = "low";

dffeas \twiddle_data[1][0][7] (
	.clk(clk),
	.d(\twiddle_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][7] .power_up = "low";

dffeas \twiddle_data[1][0][8] (
	.clk(clk),
	.d(\twiddle_data~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][8]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][8] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][8] .power_up = "low";

dffeas \twiddle_data[1][0][9] (
	.clk(clk),
	.d(\twiddle_data~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[1][0][9]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][9] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][9] .power_up = "low";

dffeas \twiddle_data[2][1][0] (
	.clk(clk),
	.d(\twiddle_data~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][0] .power_up = "low";

dffeas \twiddle_data[2][1][1] (
	.clk(clk),
	.d(\twiddle_data~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][1] .power_up = "low";

dffeas \twiddle_data[2][1][2] (
	.clk(clk),
	.d(\twiddle_data~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][2] .power_up = "low";

dffeas \twiddle_data[2][1][3] (
	.clk(clk),
	.d(\twiddle_data~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][3] .power_up = "low";

dffeas \twiddle_data[2][1][4] (
	.clk(clk),
	.d(\twiddle_data~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][4] .power_up = "low";

dffeas \twiddle_data[2][1][5] (
	.clk(clk),
	.d(\twiddle_data~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][5] .power_up = "low";

dffeas \twiddle_data[2][1][6] (
	.clk(clk),
	.d(\twiddle_data~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][6] .power_up = "low";

dffeas \twiddle_data[2][1][7] (
	.clk(clk),
	.d(\twiddle_data~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][7] .power_up = "low";

dffeas \twiddle_data[2][1][8] (
	.clk(clk),
	.d(\twiddle_data~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][8]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][8] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][8] .power_up = "low";

dffeas \twiddle_data[2][1][9] (
	.clk(clk),
	.d(\twiddle_data~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][1][9]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][9] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][9] .power_up = "low";

dffeas \twiddle_data[2][0][0] (
	.clk(clk),
	.d(\twiddle_data~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][0] .power_up = "low";

dffeas \twiddle_data[2][0][1] (
	.clk(clk),
	.d(\twiddle_data~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][1] .power_up = "low";

dffeas \twiddle_data[2][0][2] (
	.clk(clk),
	.d(\twiddle_data~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][2] .power_up = "low";

dffeas \twiddle_data[2][0][3] (
	.clk(clk),
	.d(\twiddle_data~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][3] .power_up = "low";

dffeas \twiddle_data[2][0][4] (
	.clk(clk),
	.d(\twiddle_data~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][4] .power_up = "low";

dffeas \twiddle_data[2][0][5] (
	.clk(clk),
	.d(\twiddle_data~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][5] .power_up = "low";

dffeas \twiddle_data[2][0][6] (
	.clk(clk),
	.d(\twiddle_data~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][6] .power_up = "low";

dffeas \twiddle_data[2][0][7] (
	.clk(clk),
	.d(\twiddle_data~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][7] .power_up = "low";

dffeas \twiddle_data[2][0][8] (
	.clk(clk),
	.d(\twiddle_data~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][8]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][8] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][8] .power_up = "low";

dffeas \twiddle_data[2][0][9] (
	.clk(clk),
	.d(\twiddle_data~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\twiddle_data[2][0][9]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][9] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][9] .power_up = "low";

dffeas \data_rdy_vec[12] (
	.clk(clk),
	.d(\data_rdy_vec~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[12]~q ),
	.prn(vcc));
defparam \data_rdy_vec[12] .is_wysiwyg = "true";
defparam \data_rdy_vec[12] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~14 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~14_combout ),
	.cout());
defparam \data_rdy_vec~14 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~14 .sum_lutc_input = "datac";

dffeas \p_tdl[12][2] (
	.clk(clk),
	.d(\p_tdl~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[12][2]~q ),
	.prn(vcc));
defparam \p_tdl[12][2] .is_wysiwyg = "true";
defparam \p_tdl[12][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~0 (
	.dataa(reset_n),
	.datab(\p_tdl[12][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~0_combout ),
	.cout());
defparam \p_tdl~0 .lut_mask = 16'hEEEE;
defparam \p_tdl~0 .sum_lutc_input = "datac";

dffeas \p_tdl[12][0] (
	.clk(clk),
	.d(\p_tdl~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[12][0]~q ),
	.prn(vcc));
defparam \p_tdl[12][0] .is_wysiwyg = "true";
defparam \p_tdl[12][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~1 (
	.dataa(reset_n),
	.datab(\p_tdl[12][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~1_combout ),
	.cout());
defparam \p_tdl~1 .lut_mask = 16'hEEEE;
defparam \p_tdl~1 .sum_lutc_input = "datac";

dffeas \p_tdl[12][1] (
	.clk(clk),
	.d(\p_tdl~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[12][1]~q ),
	.prn(vcc));
defparam \p_tdl[12][1] .is_wysiwyg = "true";
defparam \p_tdl[12][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~2 (
	.dataa(reset_n),
	.datab(\p_tdl[12][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~2_combout ),
	.cout());
defparam \p_tdl~2 .lut_mask = 16'hEEEE;
defparam \p_tdl~2 .sum_lutc_input = "datac";

dffeas \p_tdl[10][0] (
	.clk(clk),
	.d(\p_tdl~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[10][0]~q ),
	.prn(vcc));
defparam \p_tdl[10][0] .is_wysiwyg = "true";
defparam \p_tdl[10][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~3 (
	.dataa(reset_n),
	.datab(\p_tdl[10][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~3_combout ),
	.cout());
defparam \p_tdl~3 .lut_mask = 16'hEEEE;
defparam \p_tdl~3 .sum_lutc_input = "datac";

dffeas \p_tdl[10][2] (
	.clk(clk),
	.d(\p_tdl~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[10][2]~q ),
	.prn(vcc));
defparam \p_tdl[10][2] .is_wysiwyg = "true";
defparam \p_tdl[10][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~4 (
	.dataa(reset_n),
	.datab(\p_tdl[10][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~4_combout ),
	.cout());
defparam \p_tdl~4 .lut_mask = 16'hEEEE;
defparam \p_tdl~4 .sum_lutc_input = "datac";

dffeas \p_tdl[10][1] (
	.clk(clk),
	.d(\p_tdl~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[10][1]~q ),
	.prn(vcc));
defparam \p_tdl[10][1] .is_wysiwyg = "true";
defparam \p_tdl[10][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~5 (
	.dataa(reset_n),
	.datab(\p_tdl[10][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~5_combout ),
	.cout());
defparam \p_tdl~5 .lut_mask = 16'hEEEE;
defparam \p_tdl~5 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[3] (
	.clk(clk),
	.d(\data_rdy_vec~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[3]~q ),
	.prn(vcc));
defparam \data_rdy_vec[3] .is_wysiwyg = "true";
defparam \data_rdy_vec[3] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~15 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~15_combout ),
	.cout());
defparam \data_rdy_vec~15 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~0 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~0_combout ),
	.cout());
defparam \twiddle_data~0 .lut_mask = 16'hEEEE;
defparam \twiddle_data~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~1 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~1_combout ),
	.cout());
defparam \twiddle_data~1 .lut_mask = 16'hEEEE;
defparam \twiddle_data~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~2 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~2_combout ),
	.cout());
defparam \twiddle_data~2 .lut_mask = 16'hEEEE;
defparam \twiddle_data~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~3 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~3_combout ),
	.cout());
defparam \twiddle_data~3 .lut_mask = 16'hEEEE;
defparam \twiddle_data~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~4 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~4_combout ),
	.cout());
defparam \twiddle_data~4 .lut_mask = 16'hEEEE;
defparam \twiddle_data~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~5 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~5_combout ),
	.cout());
defparam \twiddle_data~5 .lut_mask = 16'hEEEE;
defparam \twiddle_data~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~6 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~6_combout ),
	.cout());
defparam \twiddle_data~6 .lut_mask = 16'hEEEE;
defparam \twiddle_data~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~7 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~7_combout ),
	.cout());
defparam \twiddle_data~7 .lut_mask = 16'hEEEE;
defparam \twiddle_data~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~8 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~8_combout ),
	.cout());
defparam \twiddle_data~8 .lut_mask = 16'hEEEE;
defparam \twiddle_data~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~9 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~9_combout ),
	.cout());
defparam \twiddle_data~9 .lut_mask = 16'hEEEE;
defparam \twiddle_data~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~10 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~10_combout ),
	.cout());
defparam \twiddle_data~10 .lut_mask = 16'hAAFF;
defparam \twiddle_data~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~11 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~11_combout ),
	.cout());
defparam \twiddle_data~11 .lut_mask = 16'hAAFF;
defparam \twiddle_data~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~12 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~12_combout ),
	.cout());
defparam \twiddle_data~12 .lut_mask = 16'hAAFF;
defparam \twiddle_data~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~13 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~13_combout ),
	.cout());
defparam \twiddle_data~13 .lut_mask = 16'hAAFF;
defparam \twiddle_data~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~14 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~14_combout ),
	.cout());
defparam \twiddle_data~14 .lut_mask = 16'hAAFF;
defparam \twiddle_data~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~15 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~15_combout ),
	.cout());
defparam \twiddle_data~15 .lut_mask = 16'hAAFF;
defparam \twiddle_data~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~16 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~16_combout ),
	.cout());
defparam \twiddle_data~16 .lut_mask = 16'hAAFF;
defparam \twiddle_data~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~17 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~17_combout ),
	.cout());
defparam \twiddle_data~17 .lut_mask = 16'hAAFF;
defparam \twiddle_data~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~18 (
	.dataa(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~18_combout ),
	.cout());
defparam \twiddle_data~18 .lut_mask = 16'hAAFF;
defparam \twiddle_data~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~19 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~19_combout ),
	.cout());
defparam \twiddle_data~19 .lut_mask = 16'hEEEE;
defparam \twiddle_data~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~20 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~20_combout ),
	.cout());
defparam \twiddle_data~20 .lut_mask = 16'hEEEE;
defparam \twiddle_data~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~21 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~21_combout ),
	.cout());
defparam \twiddle_data~21 .lut_mask = 16'hEEEE;
defparam \twiddle_data~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~22 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~22_combout ),
	.cout());
defparam \twiddle_data~22 .lut_mask = 16'hEEEE;
defparam \twiddle_data~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~23 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~23_combout ),
	.cout());
defparam \twiddle_data~23 .lut_mask = 16'hEEEE;
defparam \twiddle_data~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~24 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~24_combout ),
	.cout());
defparam \twiddle_data~24 .lut_mask = 16'hEEEE;
defparam \twiddle_data~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~25 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~25_combout ),
	.cout());
defparam \twiddle_data~25 .lut_mask = 16'hEEEE;
defparam \twiddle_data~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~26 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~26_combout ),
	.cout());
defparam \twiddle_data~26 .lut_mask = 16'hEEEE;
defparam \twiddle_data~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~27 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~27_combout ),
	.cout());
defparam \twiddle_data~27 .lut_mask = 16'hEEEE;
defparam \twiddle_data~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~28 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~28_combout ),
	.cout());
defparam \twiddle_data~28 .lut_mask = 16'hEEEE;
defparam \twiddle_data~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~29 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~29_combout ),
	.cout());
defparam \twiddle_data~29 .lut_mask = 16'hEEEE;
defparam \twiddle_data~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~30 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~30_combout ),
	.cout());
defparam \twiddle_data~30 .lut_mask = 16'hAAFF;
defparam \twiddle_data~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~31 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~31_combout ),
	.cout());
defparam \twiddle_data~31 .lut_mask = 16'hAAFF;
defparam \twiddle_data~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~32 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~32_combout ),
	.cout());
defparam \twiddle_data~32 .lut_mask = 16'hAAFF;
defparam \twiddle_data~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~33 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~33_combout ),
	.cout());
defparam \twiddle_data~33 .lut_mask = 16'hAAFF;
defparam \twiddle_data~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~34 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~34_combout ),
	.cout());
defparam \twiddle_data~34 .lut_mask = 16'hAAFF;
defparam \twiddle_data~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~35 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~35_combout ),
	.cout());
defparam \twiddle_data~35 .lut_mask = 16'hAAFF;
defparam \twiddle_data~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~36 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~36_combout ),
	.cout());
defparam \twiddle_data~36 .lut_mask = 16'hAAFF;
defparam \twiddle_data~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~37 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~37_combout ),
	.cout());
defparam \twiddle_data~37 .lut_mask = 16'hAAFF;
defparam \twiddle_data~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~38 (
	.dataa(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~38_combout ),
	.cout());
defparam \twiddle_data~38 .lut_mask = 16'hAAFF;
defparam \twiddle_data~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~39 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~39_combout ),
	.cout());
defparam \twiddle_data~39 .lut_mask = 16'hEEEE;
defparam \twiddle_data~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~40 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~40_combout ),
	.cout());
defparam \twiddle_data~40 .lut_mask = 16'hEEEE;
defparam \twiddle_data~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~41 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~41_combout ),
	.cout());
defparam \twiddle_data~41 .lut_mask = 16'hEEEE;
defparam \twiddle_data~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~42 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~42_combout ),
	.cout());
defparam \twiddle_data~42 .lut_mask = 16'hEEEE;
defparam \twiddle_data~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~43 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~43_combout ),
	.cout());
defparam \twiddle_data~43 .lut_mask = 16'hEEEE;
defparam \twiddle_data~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~44 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~44_combout ),
	.cout());
defparam \twiddle_data~44 .lut_mask = 16'hEEEE;
defparam \twiddle_data~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~45 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~45_combout ),
	.cout());
defparam \twiddle_data~45 .lut_mask = 16'hEEEE;
defparam \twiddle_data~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~46 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~46_combout ),
	.cout());
defparam \twiddle_data~46 .lut_mask = 16'hEEEE;
defparam \twiddle_data~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~47 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~47_combout ),
	.cout());
defparam \twiddle_data~47 .lut_mask = 16'hEEEE;
defparam \twiddle_data~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~48 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~48_combout ),
	.cout());
defparam \twiddle_data~48 .lut_mask = 16'hEEEE;
defparam \twiddle_data~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~49 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~49_combout ),
	.cout());
defparam \twiddle_data~49 .lut_mask = 16'hEEEE;
defparam \twiddle_data~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~50 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~50_combout ),
	.cout());
defparam \twiddle_data~50 .lut_mask = 16'hAAFF;
defparam \twiddle_data~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~51 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~51_combout ),
	.cout());
defparam \twiddle_data~51 .lut_mask = 16'hAAFF;
defparam \twiddle_data~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~52 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~52_combout ),
	.cout());
defparam \twiddle_data~52 .lut_mask = 16'hAAFF;
defparam \twiddle_data~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~53 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~53_combout ),
	.cout());
defparam \twiddle_data~53 .lut_mask = 16'hAAFF;
defparam \twiddle_data~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~54 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~54_combout ),
	.cout());
defparam \twiddle_data~54 .lut_mask = 16'hAAFF;
defparam \twiddle_data~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~55 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~55_combout ),
	.cout());
defparam \twiddle_data~55 .lut_mask = 16'hAAFF;
defparam \twiddle_data~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~56 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~56_combout ),
	.cout());
defparam \twiddle_data~56 .lut_mask = 16'hAAFF;
defparam \twiddle_data~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~57 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~57_combout ),
	.cout());
defparam \twiddle_data~57 .lut_mask = 16'hAAFF;
defparam \twiddle_data~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~58 (
	.dataa(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\twiddle_data~58_combout ),
	.cout());
defparam \twiddle_data~58 .lut_mask = 16'hAAFF;
defparam \twiddle_data~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twiddle_data~59 (
	.dataa(reset_n),
	.datab(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twiddle_data~59_combout ),
	.cout());
defparam \twiddle_data~59 .lut_mask = 16'hEEEE;
defparam \twiddle_data~59 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[11] (
	.clk(clk),
	.d(\data_rdy_vec~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[11]~q ),
	.prn(vcc));
defparam \data_rdy_vec[11] .is_wysiwyg = "true";
defparam \data_rdy_vec[11] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~16 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~16_combout ),
	.cout());
defparam \data_rdy_vec~16 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~6 (
	.dataa(reset_n),
	.datab(\p_tdl[11][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~6_combout ),
	.cout());
defparam \p_tdl~6 .lut_mask = 16'hEEEE;
defparam \p_tdl~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~7 (
	.dataa(reset_n),
	.datab(\p_tdl[11][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~7_combout ),
	.cout());
defparam \p_tdl~7 .lut_mask = 16'hEEEE;
defparam \p_tdl~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~8 (
	.dataa(reset_n),
	.datab(\p_tdl[11][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~8_combout ),
	.cout());
defparam \p_tdl~8 .lut_mask = 16'hEEEE;
defparam \p_tdl~8 .sum_lutc_input = "datac";

dffeas \p_tdl[9][0] (
	.clk(clk),
	.d(\p_tdl~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[9][0]~q ),
	.prn(vcc));
defparam \p_tdl[9][0] .is_wysiwyg = "true";
defparam \p_tdl[9][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~9 (
	.dataa(reset_n),
	.datab(\p_tdl[9][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~9_combout ),
	.cout());
defparam \p_tdl~9 .lut_mask = 16'hEEEE;
defparam \p_tdl~9 .sum_lutc_input = "datac";

dffeas \p_tdl[9][2] (
	.clk(clk),
	.d(\p_tdl~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[9][2]~q ),
	.prn(vcc));
defparam \p_tdl[9][2] .is_wysiwyg = "true";
defparam \p_tdl[9][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~10 (
	.dataa(reset_n),
	.datab(\p_tdl[9][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~10_combout ),
	.cout());
defparam \p_tdl~10 .lut_mask = 16'hEEEE;
defparam \p_tdl~10 .sum_lutc_input = "datac";

dffeas \p_tdl[9][1] (
	.clk(clk),
	.d(\p_tdl~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[9][1]~q ),
	.prn(vcc));
defparam \p_tdl[9][1] .is_wysiwyg = "true";
defparam \p_tdl[9][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~11 (
	.dataa(reset_n),
	.datab(\p_tdl[9][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~11_combout ),
	.cout());
defparam \p_tdl~11 .lut_mask = 16'hEEEE;
defparam \p_tdl~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_vec~17 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~17_combout ),
	.cout());
defparam \data_rdy_vec~17 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~17 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[10] (
	.clk(clk),
	.d(\data_rdy_vec~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[10]~q ),
	.prn(vcc));
defparam \data_rdy_vec[10] .is_wysiwyg = "true";
defparam \data_rdy_vec[10] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~18 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~18_combout ),
	.cout());
defparam \data_rdy_vec~18 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~18 .sum_lutc_input = "datac";

dffeas \p_tdl[8][0] (
	.clk(clk),
	.d(\p_tdl~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[8][0]~q ),
	.prn(vcc));
defparam \p_tdl[8][0] .is_wysiwyg = "true";
defparam \p_tdl[8][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~12 (
	.dataa(reset_n),
	.datab(\p_tdl[8][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~12_combout ),
	.cout());
defparam \p_tdl~12 .lut_mask = 16'hEEEE;
defparam \p_tdl~12 .sum_lutc_input = "datac";

dffeas \p_tdl[8][2] (
	.clk(clk),
	.d(\p_tdl~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[8][2]~q ),
	.prn(vcc));
defparam \p_tdl[8][2] .is_wysiwyg = "true";
defparam \p_tdl[8][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~13 (
	.dataa(reset_n),
	.datab(\p_tdl[8][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~13_combout ),
	.cout());
defparam \p_tdl~13 .lut_mask = 16'hEEEE;
defparam \p_tdl~13 .sum_lutc_input = "datac";

dffeas \p_tdl[8][1] (
	.clk(clk),
	.d(\p_tdl~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[8][1]~q ),
	.prn(vcc));
defparam \p_tdl[8][1] .is_wysiwyg = "true";
defparam \p_tdl[8][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~14 (
	.dataa(reset_n),
	.datab(\p_tdl[8][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~14_combout ),
	.cout());
defparam \p_tdl~14 .lut_mask = 16'hEEEE;
defparam \p_tdl~14 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[9] (
	.clk(clk),
	.d(\data_rdy_vec~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[9]~q ),
	.prn(vcc));
defparam \data_rdy_vec[9] .is_wysiwyg = "true";
defparam \data_rdy_vec[9] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~19 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~19_combout ),
	.cout());
defparam \data_rdy_vec~19 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~19 .sum_lutc_input = "datac";

dffeas \p_tdl[7][0] (
	.clk(clk),
	.d(\p_tdl~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[7][0]~q ),
	.prn(vcc));
defparam \p_tdl[7][0] .is_wysiwyg = "true";
defparam \p_tdl[7][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~15 (
	.dataa(reset_n),
	.datab(\p_tdl[7][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~15_combout ),
	.cout());
defparam \p_tdl~15 .lut_mask = 16'hEEEE;
defparam \p_tdl~15 .sum_lutc_input = "datac";

dffeas \p_tdl[7][2] (
	.clk(clk),
	.d(\p_tdl~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[7][2]~q ),
	.prn(vcc));
defparam \p_tdl[7][2] .is_wysiwyg = "true";
defparam \p_tdl[7][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~16 (
	.dataa(reset_n),
	.datab(\p_tdl[7][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~16_combout ),
	.cout());
defparam \p_tdl~16 .lut_mask = 16'hEEEE;
defparam \p_tdl~16 .sum_lutc_input = "datac";

dffeas \p_tdl[7][1] (
	.clk(clk),
	.d(\p_tdl~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[7][1]~q ),
	.prn(vcc));
defparam \p_tdl[7][1] .is_wysiwyg = "true";
defparam \p_tdl[7][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~17 (
	.dataa(reset_n),
	.datab(\p_tdl[7][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~17_combout ),
	.cout());
defparam \p_tdl~17 .lut_mask = 16'hEEEE;
defparam \p_tdl~17 .sum_lutc_input = "datac";

dffeas \data_rdy_vec[8] (
	.clk(clk),
	.d(\data_rdy_vec~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[8]~q ),
	.prn(vcc));
defparam \data_rdy_vec[8] .is_wysiwyg = "true";
defparam \data_rdy_vec[8] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~20 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~20_combout ),
	.cout());
defparam \data_rdy_vec~20 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~20 .sum_lutc_input = "datac";

dffeas \p_tdl[6][0] (
	.clk(clk),
	.d(\p_tdl~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[6][0]~q ),
	.prn(vcc));
defparam \p_tdl[6][0] .is_wysiwyg = "true";
defparam \p_tdl[6][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~18 (
	.dataa(reset_n),
	.datab(\p_tdl[6][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~18_combout ),
	.cout());
defparam \p_tdl~18 .lut_mask = 16'hEEEE;
defparam \p_tdl~18 .sum_lutc_input = "datac";

dffeas \p_tdl[6][2] (
	.clk(clk),
	.d(\p_tdl~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[6][2]~q ),
	.prn(vcc));
defparam \p_tdl[6][2] .is_wysiwyg = "true";
defparam \p_tdl[6][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~19 (
	.dataa(reset_n),
	.datab(\p_tdl[6][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~19_combout ),
	.cout());
defparam \p_tdl~19 .lut_mask = 16'hEEEE;
defparam \p_tdl~19 .sum_lutc_input = "datac";

dffeas \p_tdl[6][1] (
	.clk(clk),
	.d(\p_tdl~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[6][1]~q ),
	.prn(vcc));
defparam \p_tdl[6][1] .is_wysiwyg = "true";
defparam \p_tdl[6][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~20 (
	.dataa(reset_n),
	.datab(\p_tdl[6][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~20_combout ),
	.cout());
defparam \p_tdl~20 .lut_mask = 16'hEEEE;
defparam \p_tdl~20 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[4][0] (
	.clk(clk),
	.d(\sw_r_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[4][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][0] .power_up = "low";

dffeas \sw_r_tdl[4][1] (
	.clk(clk),
	.d(\sw_r_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[4][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][1] .power_up = "low";

dffeas \data_rdy_vec[7] (
	.clk(clk),
	.d(\data_rdy_vec~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[7]~q ),
	.prn(vcc));
defparam \data_rdy_vec[7] .is_wysiwyg = "true";
defparam \data_rdy_vec[7] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~21 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~21_combout ),
	.cout());
defparam \data_rdy_vec~21 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~21 .sum_lutc_input = "datac";

dffeas \p_tdl[5][0] (
	.clk(clk),
	.d(\p_tdl~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[5][0]~q ),
	.prn(vcc));
defparam \p_tdl[5][0] .is_wysiwyg = "true";
defparam \p_tdl[5][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~21 (
	.dataa(reset_n),
	.datab(\p_tdl[5][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~21_combout ),
	.cout());
defparam \p_tdl~21 .lut_mask = 16'hEEEE;
defparam \p_tdl~21 .sum_lutc_input = "datac";

dffeas \p_tdl[5][2] (
	.clk(clk),
	.d(\p_tdl~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[5][2]~q ),
	.prn(vcc));
defparam \p_tdl[5][2] .is_wysiwyg = "true";
defparam \p_tdl[5][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~22 (
	.dataa(reset_n),
	.datab(\p_tdl[5][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~22_combout ),
	.cout());
defparam \p_tdl~22 .lut_mask = 16'hEEEE;
defparam \p_tdl~22 .sum_lutc_input = "datac";

dffeas \p_tdl[5][1] (
	.clk(clk),
	.d(\p_tdl~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[5][1]~q ),
	.prn(vcc));
defparam \p_tdl[5][1] .is_wysiwyg = "true";
defparam \p_tdl[5][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~23 (
	.dataa(reset_n),
	.datab(\p_tdl[5][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~23_combout ),
	.cout());
defparam \p_tdl~23 .lut_mask = 16'hEEEE;
defparam \p_tdl~23 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[3][0] (
	.clk(clk),
	.d(\sw_r_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[3][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][0] .power_up = "low";

dffeas \sw_r_tdl[3][1] (
	.clk(clk),
	.d(\sw_r_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[3][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][1] .power_up = "low";

dffeas \data_rdy_vec[6] (
	.clk(clk),
	.d(\data_rdy_vec~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[6]~q ),
	.prn(vcc));
defparam \data_rdy_vec[6] .is_wysiwyg = "true";
defparam \data_rdy_vec[6] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~22 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~22_combout ),
	.cout());
defparam \data_rdy_vec~22 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~22 .sum_lutc_input = "datac";

dffeas \p_tdl[4][0] (
	.clk(clk),
	.d(\p_tdl~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[4][0]~q ),
	.prn(vcc));
defparam \p_tdl[4][0] .is_wysiwyg = "true";
defparam \p_tdl[4][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~24 (
	.dataa(reset_n),
	.datab(\p_tdl[4][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~24_combout ),
	.cout());
defparam \p_tdl~24 .lut_mask = 16'hEEEE;
defparam \p_tdl~24 .sum_lutc_input = "datac";

dffeas \p_tdl[4][2] (
	.clk(clk),
	.d(\p_tdl~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[4][2]~q ),
	.prn(vcc));
defparam \p_tdl[4][2] .is_wysiwyg = "true";
defparam \p_tdl[4][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~25 (
	.dataa(reset_n),
	.datab(\p_tdl[4][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~25_combout ),
	.cout());
defparam \p_tdl~25 .lut_mask = 16'hEEEE;
defparam \p_tdl~25 .sum_lutc_input = "datac";

dffeas \p_tdl[4][1] (
	.clk(clk),
	.d(\p_tdl~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[4][1]~q ),
	.prn(vcc));
defparam \p_tdl[4][1] .is_wysiwyg = "true";
defparam \p_tdl[4][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~26 (
	.dataa(reset_n),
	.datab(\p_tdl[4][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~26_combout ),
	.cout());
defparam \p_tdl~26 .lut_mask = 16'hEEEE;
defparam \p_tdl~26 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[2][0] (
	.clk(clk),
	.d(\sw_r_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[2][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][0] .power_up = "low";

dffeas \sw_r_tdl[2][1] (
	.clk(clk),
	.d(\sw_r_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[2][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][1] .power_up = "low";

dffeas \data_rdy_vec[5] (
	.clk(clk),
	.d(\data_rdy_vec~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\data_rdy_vec[5]~q ),
	.prn(vcc));
defparam \data_rdy_vec[5] .is_wysiwyg = "true";
defparam \data_rdy_vec[5] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~23 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~23_combout ),
	.cout());
defparam \data_rdy_vec~23 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~23 .sum_lutc_input = "datac";

dffeas \p_tdl[3][0] (
	.clk(clk),
	.d(\p_tdl~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[3][0]~q ),
	.prn(vcc));
defparam \p_tdl[3][0] .is_wysiwyg = "true";
defparam \p_tdl[3][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~27 (
	.dataa(reset_n),
	.datab(\p_tdl[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~27_combout ),
	.cout());
defparam \p_tdl~27 .lut_mask = 16'hEEEE;
defparam \p_tdl~27 .sum_lutc_input = "datac";

dffeas \p_tdl[3][2] (
	.clk(clk),
	.d(\p_tdl~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[3][2]~q ),
	.prn(vcc));
defparam \p_tdl[3][2] .is_wysiwyg = "true";
defparam \p_tdl[3][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~28 (
	.dataa(reset_n),
	.datab(\p_tdl[3][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~28_combout ),
	.cout());
defparam \p_tdl~28 .lut_mask = 16'hEEEE;
defparam \p_tdl~28 .sum_lutc_input = "datac";

dffeas \p_tdl[3][1] (
	.clk(clk),
	.d(\p_tdl~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[3][1]~q ),
	.prn(vcc));
defparam \p_tdl[3][1] .is_wysiwyg = "true";
defparam \p_tdl[3][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~29 (
	.dataa(reset_n),
	.datab(\p_tdl[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~29_combout ),
	.cout());
defparam \p_tdl~29 .lut_mask = 16'hEEEE;
defparam \p_tdl~29 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[1][0] (
	.clk(clk),
	.d(\sw_r_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[1][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][0] .power_up = "low";

dffeas \sw_r_tdl[1][1] (
	.clk(clk),
	.d(\sw_r_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[1][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][1] .power_up = "low";

cycloneive_lcell_comb \data_rdy_vec~24 (
	.dataa(reset_n),
	.datab(\data_rdy_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_rdy_vec~24_combout ),
	.cout());
defparam \data_rdy_vec~24 .lut_mask = 16'hEEEE;
defparam \data_rdy_vec~24 .sum_lutc_input = "datac";

dffeas \p_tdl[2][0] (
	.clk(clk),
	.d(\p_tdl~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[2][0]~q ),
	.prn(vcc));
defparam \p_tdl[2][0] .is_wysiwyg = "true";
defparam \p_tdl[2][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~30 (
	.dataa(reset_n),
	.datab(\p_tdl[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~30_combout ),
	.cout());
defparam \p_tdl~30 .lut_mask = 16'hEEEE;
defparam \p_tdl~30 .sum_lutc_input = "datac";

dffeas \p_tdl[2][2] (
	.clk(clk),
	.d(\p_tdl~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[2][2]~q ),
	.prn(vcc));
defparam \p_tdl[2][2] .is_wysiwyg = "true";
defparam \p_tdl[2][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~31 (
	.dataa(reset_n),
	.datab(\p_tdl[2][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~31_combout ),
	.cout());
defparam \p_tdl~31 .lut_mask = 16'hEEEE;
defparam \p_tdl~31 .sum_lutc_input = "datac";

dffeas \p_tdl[2][1] (
	.clk(clk),
	.d(\p_tdl~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[2][1]~q ),
	.prn(vcc));
defparam \p_tdl[2][1] .is_wysiwyg = "true";
defparam \p_tdl[2][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~32 (
	.dataa(reset_n),
	.datab(\p_tdl[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~32_combout ),
	.cout());
defparam \p_tdl~32 .lut_mask = 16'hEEEE;
defparam \p_tdl~32 .sum_lutc_input = "datac";

dffeas \sw_r_tdl[0][0] (
	.clk(clk),
	.d(\rd_adgen|sw[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[0][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][0] .power_up = "low";

dffeas \sw_r_tdl[0][1] (
	.clk(clk),
	.d(\rd_adgen|sw[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\sw_r_tdl[0][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][1] .power_up = "low";

dffeas \p_tdl[1][0] (
	.clk(clk),
	.d(\p_tdl~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[1][0]~q ),
	.prn(vcc));
defparam \p_tdl[1][0] .is_wysiwyg = "true";
defparam \p_tdl[1][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~33 (
	.dataa(reset_n),
	.datab(\p_tdl[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~33_combout ),
	.cout());
defparam \p_tdl~33 .lut_mask = 16'hEEEE;
defparam \p_tdl~33 .sum_lutc_input = "datac";

dffeas \p_tdl[1][2] (
	.clk(clk),
	.d(\p_tdl~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[1][2]~q ),
	.prn(vcc));
defparam \p_tdl[1][2] .is_wysiwyg = "true";
defparam \p_tdl[1][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~34 (
	.dataa(reset_n),
	.datab(\p_tdl[1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~34_combout ),
	.cout());
defparam \p_tdl~34 .lut_mask = 16'hEEEE;
defparam \p_tdl~34 .sum_lutc_input = "datac";

dffeas \p_tdl[1][1] (
	.clk(clk),
	.d(\p_tdl~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[1][1]~q ),
	.prn(vcc));
defparam \p_tdl[1][1] .is_wysiwyg = "true";
defparam \p_tdl[1][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~35 (
	.dataa(reset_n),
	.datab(\p_tdl[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~35_combout ),
	.cout());
defparam \p_tdl~35 .lut_mask = 16'hEEEE;
defparam \p_tdl~35 .sum_lutc_input = "datac";

dffeas \p_tdl[0][0] (
	.clk(clk),
	.d(\p_tdl~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[0][0]~q ),
	.prn(vcc));
defparam \p_tdl[0][0] .is_wysiwyg = "true";
defparam \p_tdl[0][0] .power_up = "low";

cycloneive_lcell_comb \p_tdl~36 (
	.dataa(reset_n),
	.datab(\p_tdl[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~36_combout ),
	.cout());
defparam \p_tdl~36 .lut_mask = 16'hEEEE;
defparam \p_tdl~36 .sum_lutc_input = "datac";

dffeas \p_tdl[0][2] (
	.clk(clk),
	.d(\p_tdl~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[0][2]~q ),
	.prn(vcc));
defparam \p_tdl[0][2] .is_wysiwyg = "true";
defparam \p_tdl[0][2] .power_up = "low";

cycloneive_lcell_comb \p_tdl~37 (
	.dataa(reset_n),
	.datab(\p_tdl[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~37_combout ),
	.cout());
defparam \p_tdl~37 .lut_mask = 16'hEEEE;
defparam \p_tdl~37 .sum_lutc_input = "datac";

dffeas \p_tdl[0][1] (
	.clk(clk),
	.d(\p_tdl~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\global_clock_enable~1_combout ),
	.q(\p_tdl[0][1]~q ),
	.prn(vcc));
defparam \p_tdl[0][1] .is_wysiwyg = "true";
defparam \p_tdl[0][1] .power_up = "low";

cycloneive_lcell_comb \p_tdl~38 (
	.dataa(reset_n),
	.datab(\p_tdl[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~38_combout ),
	.cout());
defparam \p_tdl~38 .lut_mask = 16'hEEEE;
defparam \p_tdl~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~39 (
	.dataa(reset_n),
	.datab(\ctrl|p[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~39_combout ),
	.cout());
defparam \p_tdl~39 .lut_mask = 16'hEEEE;
defparam \p_tdl~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~40 (
	.dataa(reset_n),
	.datab(\ctrl|p[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~40_combout ),
	.cout());
defparam \p_tdl~40 .lut_mask = 16'hEEEE;
defparam \p_tdl~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p_tdl~41 (
	.dataa(reset_n),
	.datab(\ctrl|p[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_tdl~41_combout ),
	.cout());
defparam \p_tdl~41 .lut_mask = 16'hEEEE;
defparam \p_tdl~41 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_3dp_rom (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_01,
	q_a_11,
	q_a_21,
	q_a_31,
	q_a_41,
	q_a_51,
	q_a_61,
	q_a_71,
	q_a_81,
	q_a_91,
	q_a_02,
	q_a_12,
	q_a_22,
	q_a_32,
	q_a_42,
	q_a_52,
	q_a_62,
	q_a_72,
	q_a_82,
	q_a_92,
	q_a_03,
	q_a_13,
	q_a_23,
	q_a_33,
	q_a_43,
	q_a_53,
	q_a_63,
	q_a_73,
	q_a_83,
	q_a_93,
	q_a_04,
	q_a_14,
	q_a_24,
	q_a_34,
	q_a_44,
	q_a_54,
	q_a_64,
	q_a_74,
	q_a_84,
	q_a_94,
	q_a_05,
	q_a_15,
	q_a_25,
	q_a_35,
	q_a_45,
	q_a_55,
	q_a_65,
	q_a_75,
	q_a_85,
	q_a_95,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
output 	q_a_01;
output 	q_a_11;
output 	q_a_21;
output 	q_a_31;
output 	q_a_41;
output 	q_a_51;
output 	q_a_61;
output 	q_a_71;
output 	q_a_81;
output 	q_a_91;
output 	q_a_02;
output 	q_a_12;
output 	q_a_22;
output 	q_a_32;
output 	q_a_42;
output 	q_a_52;
output 	q_a_62;
output 	q_a_72;
output 	q_a_82;
output 	q_a_92;
output 	q_a_03;
output 	q_a_13;
output 	q_a_23;
output 	q_a_33;
output 	q_a_43;
output 	q_a_53;
output 	q_a_63;
output 	q_a_73;
output 	q_a_83;
output 	q_a_93;
output 	q_a_04;
output 	q_a_14;
output 	q_a_24;
output 	q_a_34;
output 	q_a_44;
output 	q_a_54;
output 	q_a_64;
output 	q_a_74;
output 	q_a_84;
output 	q_a_94;
output 	q_a_05;
output 	q_a_15;
output 	q_a_25;
output 	q_a_35;
output 	q_a_45;
output 	q_a_55;
output 	q_a_65;
output 	q_a_75;
output 	q_a_85;
output 	q_a_95;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_twid_rom_2 \gen_M4K:cos_3n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_05),
	.q_a_1(q_a_15),
	.q_a_2(q_a_25),
	.q_a_3(q_a_35),
	.q_a_4(q_a_45),
	.q_a_5(q_a_55),
	.q_a_6(q_a_65),
	.q_a_7(q_a_75),
	.q_a_8(q_a_85),
	.q_a_9(q_a_95),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_twid_rom_1 \gen_M4K:cos_2n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_03),
	.q_a_1(q_a_13),
	.q_a_2(q_a_23),
	.q_a_3(q_a_33),
	.q_a_4(q_a_43),
	.q_a_5(q_a_53),
	.q_a_6(q_a_63),
	.q_a_7(q_a_73),
	.q_a_8(q_a_83),
	.q_a_9(q_a_93),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_twid_rom \gen_M4K:cos_1n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_01),
	.q_a_1(q_a_11),
	.q_a_2(q_a_21),
	.q_a_3(q_a_31),
	.q_a_4(q_a_41),
	.q_a_5(q_a_51),
	.q_a_6(q_a_61),
	.q_a_7(q_a_71),
	.q_a_8(q_a_81),
	.q_a_9(q_a_91),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_twid_rom_5 \gen_M4K:sin_3n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_04),
	.q_a_1(q_a_14),
	.q_a_2(q_a_24),
	.q_a_3(q_a_34),
	.q_a_4(q_a_44),
	.q_a_5(q_a_54),
	.q_a_6(q_a_64),
	.q_a_7(q_a_74),
	.q_a_8(q_a_84),
	.q_a_9(q_a_94),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_twid_rom_4 \gen_M4K:sin_2n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_02),
	.q_a_1(q_a_12),
	.q_a_2(q_a_22),
	.q_a_3(q_a_32),
	.q_a_4(q_a_42),
	.q_a_5(q_a_52),
	.q_a_6(q_a_62),
	.q_a_7(q_a_72),
	.q_a_8(q_a_82),
	.q_a_9(q_a_92),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_twid_rom_3 \gen_M4K:sin_1n (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_twid_rom (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_1 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_1 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_snt3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_snt3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'hB54AB552AAAAAAAA54AD2DB64CCCE38F03FFFE078E7326D295554A5B3731E0FF;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'hC673399CCCCCCCCC993649249696B52A55555552A5296DB64CCCC638F0F01FFF;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'h52D694B5A5A5A5A5B492DB6DB24D9366CCCCCCCE6318E38E3C3C3E07F00FFFFF;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h31CE738C639C639C738E38E38E3C70E1C3C3C3C1E0F81F81FC03FE000FFFFFFF;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h0FC1F07C1F83E07C0F81F81F81FC0FE03FC03FC01FF8007FFC0001FFFFFFFFFF;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'h003FF003FF801FFC007FF8007FFC001FFFC0003FFFF8000003FFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'h00000FFFFF800003FFFFF8000003FFFFFFC000000007FFFFFFFFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'h00000000007FFFFFFFFFF80000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_1n1024cos.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_snt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule

module fftsign_twid_rom_1 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom_1 \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom_1 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_2 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_2 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_tnt3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_tnt3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'hE35D63FC69698FF192AAD98E00007C3C787C0000E336AA931FE32D2C7F8D758F;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'h1F3B2956B271F00F8E664B5AAAAAA956AD56AAAA56926670FFFC31B6AAA4CC7F;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'h00F8E732692B55552B4B6D9333333198CE67333364DB4B5AAAAA94926663C3FF;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h0007E0F1E718CCCC9926DB4969696B4A5AD29696D24926C999998C71E1E03FFF;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h00001FF01F07C3C3871E38C718E718C639CE718E31C71E3878787C0FE01FFFFF;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'h0000000FFF003FC07F01F83F07E0F83E07C1F07E0FC0FE07F807FC001FFFFFFF;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'h0000000000FFFFC000FFF800FFE007FE003FF001FFC001FFF80003FFFFFFFFFF;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'h000000000000003FFFFFF800001FFFFE00000FFFFFC0000007FFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'h0000000000000000000007FFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_2n1024cos.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_tnt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000;

endmodule

module fftsign_twid_rom_2 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom_2 \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom_2 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_3 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_unt3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_unt3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'hC92AACC0654FCA8C5619BE57E53F6CF9ACFF92AA5936DAAA63C6A9F9583519A7;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'h924CCF001CDA930C32ADC1CD49C0E5AD30FF8E66CB6DB6661FF8CD54C7C6549F;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'hE38F0FFFFC39B6A6A4CE003CDB554931C0FF81E1C71C71E1FFFF0E669552CC7F;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h56A55AAAA952DB3738F00003C7332494AA552AB56A56A54AAAAAA52DB331C3FF;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h9B366CCCCE631C383F0000003F0F1C7399CC999326CD93266666631C70F03FFF;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'hE3C78F0F0F83E03FC000000000FF03F0783C7870E1C38F1E1E1E1F03F00FFFFF;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'hFC07F00FF003FFC0000000000000FFF007FC07F01FC07F01FE01FF000FFFFFFF;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'hFFF8000FFFFC0000000000000000000FFFFC000FFFC000FFFE0000FFFFFFFFFF;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'hFFFFFFF00000000000000000000000000003FFFFFFC0000001FFFFFFFFFFFFFF;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_3n1024cos.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_unt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000;

endmodule

module fftsign_twid_rom_3 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom_3 \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom_3 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_4 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_4 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_1ot3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_1ot3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'hFE0F19D9B4A5555296C99CE3C0FFFF81E38E6664DB696A54AAAAAAAA955AA55A;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'hFFF01E1E38C66664DB6D294A95555554A95AD2D24924D9326666666673399CC6;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'hFFFFE01FC0F87878E38E318CE6666666CD93649B6DB6925B4B4B4B4B5A52D694;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'hFFFFFFE000FF807F03F03E0F078787870E1C78E38E38E39C738C738C639CE718;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'hFFFFFFFFFF00007FFC003FF007F807F80FE07F03F03F03E07C0F83F07C1F07E0;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'hFFFFFFFFFFFFFF8000003FFFF80007FFF0007FFC003FFC007FF003FF801FF800;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFC000000007FFFFFF8000003FFFFF800003FFFFE00000;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000003FFFFFFFFFFC0000000000;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_1n1024sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_1ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule

module fftsign_twid_rom_4 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom_4 \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom_4 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_5 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_5 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_2ot3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_2ot3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'h787C0000E336AA931FE32D2C7F8D758FE35D63FC69698FF192AAD98E00007C3C;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'hAD56AAAA56926670FFFC31B6AAA4CC7FFC664AAADB187FFE1CCC92D4AAAAD56A;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'hCE67333364DB4B5AAAAA94926663C3FFFF878CCC9252AAAAB5A5B64D9999CCE6;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h5AD29696D24926C999998C71E1E03FFFFFF80F0F1C63333326C92496D2D296B4;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h39CE718E31C71E3878787C0FE01FFFFFFFFFF00FE07C3C3C38F1C718E31CE738;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'h07C1F07E0FC0FE07F807FC001FFFFFFFFFFFFFF0007FC03FC0FE07E0FC1F07C0;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'h003FF001FFC001FFF80003FFFFFFFFFFFFFFFFFFFF80003FFF0007FF001FF800;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'h00000FFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFE00000;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'h00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_2n1024sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_2ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule

module fftsign_twid_rom_5 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_single_port_rom_5 \gen_auto:rom_component (
	.ram_block3a0(ram_block3a0),
	.ram_block3a1(ram_block3a1),
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.ram_block3a01(ram_block3a01),
	.ram_block3a11(ram_block3a11),
	.ram_block3a2(ram_block3a2),
	.ram_block3a3(ram_block3a3),
	.ram_block3a4(ram_block3a4),
	.ram_block3a5(ram_block3a5),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module fftsign_altera_fft_single_port_rom_5 (
	ram_block3a0,
	ram_block3a1,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	ram_block3a01,
	ram_block3a11,
	ram_block3a2,
	ram_block3a3,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block3a0;
input 	ram_block3a1;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
input 	ram_block3a01;
input 	ram_block3a11;
input 	ram_block3a2;
input 	ram_block3a3;
input 	ram_block3a4;
input 	ram_block3a5;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_6 \old_ram_gen:old_ram_component (
	.address_a({ram_block3a1,ram_block3a0,ram_block3a5,ram_block3a4,ram_block3a3,ram_block3a2,ram_block3a11,ram_block3a01}),
	.q_a({q_a_unconnected_wire_19,q_a_unconnected_wire_18,q_a_unconnected_wire_17,q_a_unconnected_wire_16,q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,
q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module fftsign_altsyncram_6 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[19:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_3ot3 auto_generated(
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.q_a({q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_3ot3 (
	address_a,
	q_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[7:0] address_a;
output 	[9:0] q_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 256'hCB3158353F2AC78CAAB6D934AA93FE6B3E6DF94FD4FB30D462A7E54C066AA926;

cycloneive_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 256'h39659FF36A4CF87C666DB492667000725523FE6AB3FC5A4C0335533C078CCDB4;

cycloneive_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 256'h07134AA5B38F0003E1E38C71E1F0007C664AAAD98FFF9C96A96CCF03F80F0E38;

cycloneive_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 256'h00F0C66C96A555554AB5295AB55AAAD52D2666387FFFE0E732496A55555AA56A;

cycloneive_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 256'h000FC1E38E633333266C9B366CC999CCE31E1E07FFFFFF07C38E73999993364C;

cycloneive_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 256'h00003FE07E1F0F0F1E1C78F1E3C787C3E0FE01FFFFFFFFF803F07C1E1E1C3870;

cycloneive_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 256'h0000001FFE00FF00FE03F80FE03F803FE001FFFFFFFFFFFFFC007FE01FE03F80;

cycloneive_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 256'h0000000001FFFF0001FFF8001FFF80001FFFFFFFFFFFFFFFFFFF80001FFFC000;

cycloneive_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = 256'h00000000000000FFFFFFF80000007FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;

cycloneive_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "fftsign_fft_ii_0_3n1024sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_3ot3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = 256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000;

endmodule

module fftsign_asj_fft_4dp_ram (
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_1,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_19,
	q_b_191,
	q_b_192,
	q_b_193,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_18,
	q_b_181,
	q_b_182,
	q_b_183,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_17,
	q_b_171,
	q_b_172,
	q_b_173,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_16,
	q_b_161,
	q_b_162,
	q_b_163,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_154,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_144,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	global_clock_enable,
	wren_a_3,
	a_ram_data_in_bus_12,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_18,
	wraddress_a_bus_3,
	wraddress_a_bus_20,
	wraddress_a_bus_5,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_18,
	rdaddress_a_bus_3,
	rdaddress_a_bus_20,
	rdaddress_a_bus_5,
	rdaddress_a_bus_22,
	rdaddress_a_bus_7,
	wren_a_0,
	a_ram_data_in_bus_72,
	wraddress_a_bus_24,
	wraddress_a_bus_25,
	wraddress_a_bus_10,
	wraddress_a_bus_27,
	wraddress_a_bus_12,
	wraddress_a_bus_29,
	rdaddress_a_bus_24,
	rdaddress_a_bus_25,
	rdaddress_a_bus_10,
	rdaddress_a_bus_27,
	rdaddress_a_bus_12,
	rdaddress_a_bus_29,
	rdaddress_a_bus_14,
	rdaddress_a_bus_31,
	wren_a_1,
	a_ram_data_in_bus_52,
	wraddress_a_bus_17,
	wraddress_a_bus_19,
	wraddress_a_bus_21,
	rdaddress_a_bus_17,
	rdaddress_a_bus_19,
	rdaddress_a_bus_21,
	rdaddress_a_bus_23,
	wren_a_2,
	a_ram_data_in_bus_32,
	wraddress_a_bus_9,
	wraddress_a_bus_11,
	wraddress_a_bus_13,
	rdaddress_a_bus_9,
	rdaddress_a_bus_11,
	rdaddress_a_bus_13,
	rdaddress_a_bus_15,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_71,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_70,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_79,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_69,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_78,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_68,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_77,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_67,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_76,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_66,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_75,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_65,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_74,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_64,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_73,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_23,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_1;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
output 	q_b_19;
output 	q_b_191;
output 	q_b_192;
output 	q_b_193;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_18;
output 	q_b_181;
output 	q_b_182;
output 	q_b_183;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_17;
output 	q_b_171;
output 	q_b_172;
output 	q_b_173;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_16;
output 	q_b_161;
output 	q_b_162;
output 	q_b_163;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_154;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_144;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_134;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
input 	global_clock_enable;
input 	wren_a_3;
input 	a_ram_data_in_bus_12;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_20;
input 	wraddress_a_bus_5;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_20;
input 	rdaddress_a_bus_5;
input 	rdaddress_a_bus_22;
input 	rdaddress_a_bus_7;
input 	wren_a_0;
input 	a_ram_data_in_bus_72;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_25;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_27;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_29;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_25;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_27;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_29;
input 	rdaddress_a_bus_14;
input 	rdaddress_a_bus_31;
input 	wren_a_1;
input 	a_ram_data_in_bus_52;
input 	wraddress_a_bus_17;
input 	wraddress_a_bus_19;
input 	wraddress_a_bus_21;
input 	rdaddress_a_bus_17;
input 	rdaddress_a_bus_19;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_23;
input 	wren_a_2;
input 	a_ram_data_in_bus_32;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_13;
input 	rdaddress_a_bus_15;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_62;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_71;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_70;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_79;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_69;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_78;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_68;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_77;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_67;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_76;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_66;
input 	a_ram_data_in_bus_46;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_75;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_65;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_74;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_64;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_73;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_23;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_asj_fft_data_ram_3 \gen_rams:3:dat_A (
	.q_b_12(q_b_12),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_1(q_b_1),
	.q_b_10(q_b_10),
	.q_b_0(q_b_0),
	.q_b_19(q_b_19),
	.q_b_9(q_b_9),
	.q_b_18(q_b_18),
	.q_b_8(q_b_8),
	.q_b_17(q_b_17),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_6(q_b_6),
	.q_b_15(q_b_151),
	.q_b_5(q_b_5),
	.q_b_14(q_b_141),
	.q_b_4(q_b_4),
	.q_b_13(q_b_131),
	.q_b_3(q_b_3),
	.global_clock_enable(global_clock_enable),
	.wren_a_3(wren_a_3),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.wraddress_a_bus_3(wraddress_a_bus_3),
	.wraddress_a_bus_20(wraddress_a_bus_20),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.rdaddress_a_bus_3(rdaddress_a_bus_3),
	.rdaddress_a_bus_20(rdaddress_a_bus_20),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.rdaddress_a_bus_22(rdaddress_a_bus_22),
	.rdaddress_a_bus_7(rdaddress_a_bus_7),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.clk(clk));

fftsign_asj_fft_data_ram_2 \gen_rams:2:dat_A (
	.q_b_12(q_b_123),
	.q_b_2(q_b_23),
	.q_b_11(q_b_113),
	.q_b_1(q_b_15),
	.q_b_10(q_b_103),
	.q_b_0(q_b_03),
	.q_b_19(q_b_193),
	.q_b_9(q_b_93),
	.q_b_18(q_b_183),
	.q_b_8(q_b_83),
	.q_b_17(q_b_173),
	.q_b_7(q_b_73),
	.q_b_16(q_b_163),
	.q_b_6(q_b_63),
	.q_b_15(q_b_154),
	.q_b_5(q_b_53),
	.q_b_14(q_b_144),
	.q_b_4(q_b_43),
	.q_b_13(q_b_134),
	.q_b_3(q_b_33),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.wraddress_a_bus_24(wraddress_a_bus_24),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.rdaddress_a_bus_24(rdaddress_a_bus_24),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_14(rdaddress_a_bus_14),
	.wren_a_2(wren_a_2),
	.a_ram_data_in_bus_32(a_ram_data_in_bus_32),
	.wraddress_a_bus_9(wraddress_a_bus_9),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_9(rdaddress_a_bus_9),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.rdaddress_a_bus_15(rdaddress_a_bus_15),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_39(a_ram_data_in_bus_39),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_38(a_ram_data_in_bus_38),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_37(a_ram_data_in_bus_37),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_36(a_ram_data_in_bus_36),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.a_ram_data_in_bus_35(a_ram_data_in_bus_35),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_34(a_ram_data_in_bus_34),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_33(a_ram_data_in_bus_33),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.clk(clk));

fftsign_asj_fft_data_ram_1 \gen_rams:1:dat_A (
	.q_b_12(q_b_122),
	.q_b_2(q_b_22),
	.q_b_11(q_b_112),
	.q_b_1(q_b_14),
	.q_b_10(q_b_102),
	.q_b_0(q_b_02),
	.q_b_19(q_b_192),
	.q_b_9(q_b_92),
	.q_b_18(q_b_182),
	.q_b_8(q_b_82),
	.q_b_17(q_b_172),
	.q_b_7(q_b_72),
	.q_b_16(q_b_162),
	.q_b_6(q_b_62),
	.q_b_15(q_b_153),
	.q_b_5(q_b_52),
	.q_b_14(q_b_143),
	.q_b_4(q_b_42),
	.q_b_13(q_b_133),
	.q_b_3(q_b_32),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.wraddress_a_bus_20(wraddress_a_bus_20),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.rdaddress_a_bus_20(rdaddress_a_bus_20),
	.rdaddress_a_bus_22(rdaddress_a_bus_22),
	.wren_a_1(wren_a_1),
	.a_ram_data_in_bus_52(a_ram_data_in_bus_52),
	.wraddress_a_bus_17(wraddress_a_bus_17),
	.wraddress_a_bus_19(wraddress_a_bus_19),
	.wraddress_a_bus_21(wraddress_a_bus_21),
	.rdaddress_a_bus_17(rdaddress_a_bus_17),
	.rdaddress_a_bus_19(rdaddress_a_bus_19),
	.rdaddress_a_bus_21(rdaddress_a_bus_21),
	.rdaddress_a_bus_23(rdaddress_a_bus_23),
	.a_ram_data_in_bus_42(a_ram_data_in_bus_42),
	.a_ram_data_in_bus_51(a_ram_data_in_bus_51),
	.a_ram_data_in_bus_41(a_ram_data_in_bus_41),
	.a_ram_data_in_bus_50(a_ram_data_in_bus_50),
	.a_ram_data_in_bus_40(a_ram_data_in_bus_40),
	.a_ram_data_in_bus_59(a_ram_data_in_bus_59),
	.a_ram_data_in_bus_49(a_ram_data_in_bus_49),
	.a_ram_data_in_bus_58(a_ram_data_in_bus_58),
	.a_ram_data_in_bus_48(a_ram_data_in_bus_48),
	.a_ram_data_in_bus_57(a_ram_data_in_bus_57),
	.a_ram_data_in_bus_47(a_ram_data_in_bus_47),
	.a_ram_data_in_bus_56(a_ram_data_in_bus_56),
	.a_ram_data_in_bus_46(a_ram_data_in_bus_46),
	.a_ram_data_in_bus_55(a_ram_data_in_bus_55),
	.a_ram_data_in_bus_45(a_ram_data_in_bus_45),
	.a_ram_data_in_bus_54(a_ram_data_in_bus_54),
	.a_ram_data_in_bus_44(a_ram_data_in_bus_44),
	.a_ram_data_in_bus_53(a_ram_data_in_bus_53),
	.a_ram_data_in_bus_43(a_ram_data_in_bus_43),
	.clk(clk));

fftsign_asj_fft_data_ram \gen_rams:0:dat_A (
	.q_b_12(q_b_121),
	.q_b_2(q_b_21),
	.q_b_11(q_b_111),
	.q_b_1(q_b_13),
	.q_b_10(q_b_101),
	.q_b_0(q_b_01),
	.q_b_19(q_b_191),
	.q_b_9(q_b_91),
	.q_b_18(q_b_181),
	.q_b_8(q_b_81),
	.q_b_17(q_b_171),
	.q_b_7(q_b_71),
	.q_b_16(q_b_161),
	.q_b_6(q_b_61),
	.q_b_15(q_b_152),
	.q_b_5(q_b_51),
	.q_b_14(q_b_142),
	.q_b_4(q_b_41),
	.q_b_13(q_b_132),
	.q_b_3(q_b_31),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.wren_a_0(wren_a_0),
	.a_ram_data_in_bus_72(a_ram_data_in_bus_72),
	.wraddress_a_bus_24(wraddress_a_bus_24),
	.wraddress_a_bus_25(wraddress_a_bus_25),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_27(wraddress_a_bus_27),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.wraddress_a_bus_29(wraddress_a_bus_29),
	.rdaddress_a_bus_24(rdaddress_a_bus_24),
	.rdaddress_a_bus_25(rdaddress_a_bus_25),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_27(rdaddress_a_bus_27),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_29(rdaddress_a_bus_29),
	.rdaddress_a_bus_14(rdaddress_a_bus_14),
	.rdaddress_a_bus_31(rdaddress_a_bus_31),
	.a_ram_data_in_bus_62(a_ram_data_in_bus_62),
	.a_ram_data_in_bus_71(a_ram_data_in_bus_71),
	.a_ram_data_in_bus_61(a_ram_data_in_bus_61),
	.a_ram_data_in_bus_70(a_ram_data_in_bus_70),
	.a_ram_data_in_bus_60(a_ram_data_in_bus_60),
	.a_ram_data_in_bus_79(a_ram_data_in_bus_79),
	.a_ram_data_in_bus_69(a_ram_data_in_bus_69),
	.a_ram_data_in_bus_78(a_ram_data_in_bus_78),
	.a_ram_data_in_bus_68(a_ram_data_in_bus_68),
	.a_ram_data_in_bus_77(a_ram_data_in_bus_77),
	.a_ram_data_in_bus_67(a_ram_data_in_bus_67),
	.a_ram_data_in_bus_76(a_ram_data_in_bus_76),
	.a_ram_data_in_bus_66(a_ram_data_in_bus_66),
	.a_ram_data_in_bus_75(a_ram_data_in_bus_75),
	.a_ram_data_in_bus_65(a_ram_data_in_bus_65),
	.a_ram_data_in_bus_74(a_ram_data_in_bus_74),
	.a_ram_data_in_bus_64(a_ram_data_in_bus_64),
	.a_ram_data_in_bus_73(a_ram_data_in_bus_73),
	.a_ram_data_in_bus_63(a_ram_data_in_bus_63),
	.clk(clk));

endmodule

module fftsign_asj_fft_data_ram (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	wren_a_0,
	a_ram_data_in_bus_72,
	wraddress_a_bus_24,
	wraddress_a_bus_25,
	wraddress_a_bus_10,
	wraddress_a_bus_27,
	wraddress_a_bus_12,
	wraddress_a_bus_29,
	rdaddress_a_bus_24,
	rdaddress_a_bus_25,
	rdaddress_a_bus_10,
	rdaddress_a_bus_27,
	rdaddress_a_bus_12,
	rdaddress_a_bus_29,
	rdaddress_a_bus_14,
	rdaddress_a_bus_31,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_71,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_70,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_79,
	a_ram_data_in_bus_69,
	a_ram_data_in_bus_78,
	a_ram_data_in_bus_68,
	a_ram_data_in_bus_77,
	a_ram_data_in_bus_67,
	a_ram_data_in_bus_76,
	a_ram_data_in_bus_66,
	a_ram_data_in_bus_75,
	a_ram_data_in_bus_65,
	a_ram_data_in_bus_74,
	a_ram_data_in_bus_64,
	a_ram_data_in_bus_73,
	a_ram_data_in_bus_63,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	wren_a_0;
input 	a_ram_data_in_bus_72;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_25;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_27;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_29;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_25;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_27;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_29;
input 	rdaddress_a_bus_14;
input 	rdaddress_a_bus_31;
input 	a_ram_data_in_bus_62;
input 	a_ram_data_in_bus_71;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_70;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_79;
input 	a_ram_data_in_bus_69;
input 	a_ram_data_in_bus_78;
input 	a_ram_data_in_bus_68;
input 	a_ram_data_in_bus_77;
input 	a_ram_data_in_bus_67;
input 	a_ram_data_in_bus_76;
input 	a_ram_data_in_bus_66;
input 	a_ram_data_in_bus_75;
input 	a_ram_data_in_bus_65;
input 	a_ram_data_in_bus_74;
input 	a_ram_data_in_bus_64;
input 	a_ram_data_in_bus_73;
input 	a_ram_data_in_bus_63;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_dual_port_ram \gen_M4K:ram_component (
	.q_b_12(q_b_12),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_1(q_b_1),
	.q_b_10(q_b_10),
	.q_b_0(q_b_0),
	.q_b_19(q_b_19),
	.q_b_9(q_b_9),
	.q_b_18(q_b_18),
	.q_b_8(q_b_8),
	.q_b_17(q_b_17),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_3(q_b_3),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.wren_a_0(wren_a_0),
	.a_ram_data_in_bus_72(a_ram_data_in_bus_72),
	.wraddress_a_bus_24(wraddress_a_bus_24),
	.wraddress_a_bus_25(wraddress_a_bus_25),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_27(wraddress_a_bus_27),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.wraddress_a_bus_29(wraddress_a_bus_29),
	.rdaddress_a_bus_24(rdaddress_a_bus_24),
	.rdaddress_a_bus_25(rdaddress_a_bus_25),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_27(rdaddress_a_bus_27),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_29(rdaddress_a_bus_29),
	.rdaddress_a_bus_14(rdaddress_a_bus_14),
	.rdaddress_a_bus_31(rdaddress_a_bus_31),
	.a_ram_data_in_bus_62(a_ram_data_in_bus_62),
	.a_ram_data_in_bus_71(a_ram_data_in_bus_71),
	.a_ram_data_in_bus_61(a_ram_data_in_bus_61),
	.a_ram_data_in_bus_70(a_ram_data_in_bus_70),
	.a_ram_data_in_bus_60(a_ram_data_in_bus_60),
	.a_ram_data_in_bus_79(a_ram_data_in_bus_79),
	.a_ram_data_in_bus_69(a_ram_data_in_bus_69),
	.a_ram_data_in_bus_78(a_ram_data_in_bus_78),
	.a_ram_data_in_bus_68(a_ram_data_in_bus_68),
	.a_ram_data_in_bus_77(a_ram_data_in_bus_77),
	.a_ram_data_in_bus_67(a_ram_data_in_bus_67),
	.a_ram_data_in_bus_76(a_ram_data_in_bus_76),
	.a_ram_data_in_bus_66(a_ram_data_in_bus_66),
	.a_ram_data_in_bus_75(a_ram_data_in_bus_75),
	.a_ram_data_in_bus_65(a_ram_data_in_bus_65),
	.a_ram_data_in_bus_74(a_ram_data_in_bus_74),
	.a_ram_data_in_bus_64(a_ram_data_in_bus_64),
	.a_ram_data_in_bus_73(a_ram_data_in_bus_73),
	.a_ram_data_in_bus_63(a_ram_data_in_bus_63),
	.clk(clk));

endmodule

module fftsign_altera_fft_dual_port_ram (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	wren_a_0,
	a_ram_data_in_bus_72,
	wraddress_a_bus_24,
	wraddress_a_bus_25,
	wraddress_a_bus_10,
	wraddress_a_bus_27,
	wraddress_a_bus_12,
	wraddress_a_bus_29,
	rdaddress_a_bus_24,
	rdaddress_a_bus_25,
	rdaddress_a_bus_10,
	rdaddress_a_bus_27,
	rdaddress_a_bus_12,
	rdaddress_a_bus_29,
	rdaddress_a_bus_14,
	rdaddress_a_bus_31,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_71,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_70,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_79,
	a_ram_data_in_bus_69,
	a_ram_data_in_bus_78,
	a_ram_data_in_bus_68,
	a_ram_data_in_bus_77,
	a_ram_data_in_bus_67,
	a_ram_data_in_bus_76,
	a_ram_data_in_bus_66,
	a_ram_data_in_bus_75,
	a_ram_data_in_bus_65,
	a_ram_data_in_bus_74,
	a_ram_data_in_bus_64,
	a_ram_data_in_bus_73,
	a_ram_data_in_bus_63,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	wren_a_0;
input 	a_ram_data_in_bus_72;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_25;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_27;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_29;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_25;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_27;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_29;
input 	rdaddress_a_bus_14;
input 	rdaddress_a_bus_31;
input 	a_ram_data_in_bus_62;
input 	a_ram_data_in_bus_71;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_70;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_79;
input 	a_ram_data_in_bus_69;
input 	a_ram_data_in_bus_78;
input 	a_ram_data_in_bus_68;
input 	a_ram_data_in_bus_77;
input 	a_ram_data_in_bus_67;
input 	a_ram_data_in_bus_76;
input 	a_ram_data_in_bus_66;
input 	a_ram_data_in_bus_75;
input 	a_ram_data_in_bus_65;
input 	a_ram_data_in_bus_74;
input 	a_ram_data_in_bus_64;
input 	a_ram_data_in_bus_73;
input 	a_ram_data_in_bus_63;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_7 \old_ram_gen:old_ram_component (
	.q_b({q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_15,wraddress_a_bus_14,wraddress_a_bus_29,wraddress_a_bus_12,wraddress_a_bus_27,wraddress_a_bus_10,wraddress_a_bus_25,wraddress_a_bus_24}),
	.wren_a(wren_a_0),
	.data_a({a_ram_data_in_bus_79,a_ram_data_in_bus_78,a_ram_data_in_bus_77,a_ram_data_in_bus_76,a_ram_data_in_bus_75,a_ram_data_in_bus_74,a_ram_data_in_bus_73,a_ram_data_in_bus_72,a_ram_data_in_bus_71,a_ram_data_in_bus_70,a_ram_data_in_bus_69,a_ram_data_in_bus_68,
a_ram_data_in_bus_67,a_ram_data_in_bus_66,a_ram_data_in_bus_65,a_ram_data_in_bus_64,a_ram_data_in_bus_63,a_ram_data_in_bus_62,a_ram_data_in_bus_61,a_ram_data_in_bus_60}),
	.address_b({rdaddress_a_bus_31,rdaddress_a_bus_14,rdaddress_a_bus_29,rdaddress_a_bus_12,rdaddress_a_bus_27,rdaddress_a_bus_10,rdaddress_a_bus_25,rdaddress_a_bus_24}),
	.clock0(clk));

endmodule

module fftsign_altsyncram_7 (
	q_b,
	clocken0,
	address_a,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	wren_a;
input 	[19:0] data_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_d0q3 auto_generated(
	.q_b({q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clocken0(clocken0),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.data_a({data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_d0q3 (
	q_b,
	clocken0,
	address_a,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	wren_a;
input 	[19:0] data_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 20;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 20;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 20;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 20;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 20;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 20;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 20;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 20;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 20;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 20;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 20;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 20;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 20;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "clear0";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "clear0";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 20;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 20;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 20;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 20;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "clear0";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "clear0";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 20;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 20;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 20;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 20;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "clear0";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "clear0";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 20;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 20;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 20;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 20;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "clear0";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "clear0";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 20;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 20;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 20;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 20;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 20;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 20;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 20;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 20;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 20;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 20;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 20;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 20;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 20;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 20;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 20;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module fftsign_asj_fft_data_ram_1 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_0,
	wraddress_a_bus_18,
	wraddress_a_bus_20,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_18,
	rdaddress_a_bus_20,
	rdaddress_a_bus_22,
	wren_a_1,
	a_ram_data_in_bus_52,
	wraddress_a_bus_17,
	wraddress_a_bus_19,
	wraddress_a_bus_21,
	rdaddress_a_bus_17,
	rdaddress_a_bus_19,
	rdaddress_a_bus_21,
	rdaddress_a_bus_23,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_43,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_20;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_20;
input 	rdaddress_a_bus_22;
input 	wren_a_1;
input 	a_ram_data_in_bus_52;
input 	wraddress_a_bus_17;
input 	wraddress_a_bus_19;
input 	wraddress_a_bus_21;
input 	rdaddress_a_bus_17;
input 	rdaddress_a_bus_19;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_23;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_46;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_43;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_dual_port_ram_1 \gen_M4K:ram_component (
	.q_b_12(q_b_12),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_1(q_b_1),
	.q_b_10(q_b_10),
	.q_b_0(q_b_0),
	.q_b_19(q_b_19),
	.q_b_9(q_b_9),
	.q_b_18(q_b_18),
	.q_b_8(q_b_8),
	.q_b_17(q_b_17),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_3(q_b_3),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.wraddress_a_bus_20(wraddress_a_bus_20),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.rdaddress_a_bus_20(rdaddress_a_bus_20),
	.rdaddress_a_bus_22(rdaddress_a_bus_22),
	.wren_a_1(wren_a_1),
	.a_ram_data_in_bus_52(a_ram_data_in_bus_52),
	.wraddress_a_bus_17(wraddress_a_bus_17),
	.wraddress_a_bus_19(wraddress_a_bus_19),
	.wraddress_a_bus_21(wraddress_a_bus_21),
	.rdaddress_a_bus_17(rdaddress_a_bus_17),
	.rdaddress_a_bus_19(rdaddress_a_bus_19),
	.rdaddress_a_bus_21(rdaddress_a_bus_21),
	.rdaddress_a_bus_23(rdaddress_a_bus_23),
	.a_ram_data_in_bus_42(a_ram_data_in_bus_42),
	.a_ram_data_in_bus_51(a_ram_data_in_bus_51),
	.a_ram_data_in_bus_41(a_ram_data_in_bus_41),
	.a_ram_data_in_bus_50(a_ram_data_in_bus_50),
	.a_ram_data_in_bus_40(a_ram_data_in_bus_40),
	.a_ram_data_in_bus_59(a_ram_data_in_bus_59),
	.a_ram_data_in_bus_49(a_ram_data_in_bus_49),
	.a_ram_data_in_bus_58(a_ram_data_in_bus_58),
	.a_ram_data_in_bus_48(a_ram_data_in_bus_48),
	.a_ram_data_in_bus_57(a_ram_data_in_bus_57),
	.a_ram_data_in_bus_47(a_ram_data_in_bus_47),
	.a_ram_data_in_bus_56(a_ram_data_in_bus_56),
	.a_ram_data_in_bus_46(a_ram_data_in_bus_46),
	.a_ram_data_in_bus_55(a_ram_data_in_bus_55),
	.a_ram_data_in_bus_45(a_ram_data_in_bus_45),
	.a_ram_data_in_bus_54(a_ram_data_in_bus_54),
	.a_ram_data_in_bus_44(a_ram_data_in_bus_44),
	.a_ram_data_in_bus_53(a_ram_data_in_bus_53),
	.a_ram_data_in_bus_43(a_ram_data_in_bus_43),
	.clk(clk));

endmodule

module fftsign_altera_fft_dual_port_ram_1 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_0,
	wraddress_a_bus_18,
	wraddress_a_bus_20,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_18,
	rdaddress_a_bus_20,
	rdaddress_a_bus_22,
	wren_a_1,
	a_ram_data_in_bus_52,
	wraddress_a_bus_17,
	wraddress_a_bus_19,
	wraddress_a_bus_21,
	rdaddress_a_bus_17,
	rdaddress_a_bus_19,
	rdaddress_a_bus_21,
	rdaddress_a_bus_23,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_43,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_20;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_20;
input 	rdaddress_a_bus_22;
input 	wren_a_1;
input 	a_ram_data_in_bus_52;
input 	wraddress_a_bus_17;
input 	wraddress_a_bus_19;
input 	wraddress_a_bus_21;
input 	rdaddress_a_bus_17;
input 	rdaddress_a_bus_19;
input 	rdaddress_a_bus_21;
input 	rdaddress_a_bus_23;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_46;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_43;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_8 \old_ram_gen:old_ram_component (
	.q_b({q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_15,wraddress_a_bus_14,wraddress_a_bus_21,wraddress_a_bus_20,wraddress_a_bus_19,wraddress_a_bus_18,wraddress_a_bus_17,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_23,rdaddress_a_bus_22,rdaddress_a_bus_21,rdaddress_a_bus_20,rdaddress_a_bus_19,rdaddress_a_bus_18,rdaddress_a_bus_17,rdaddress_a_bus_0}),
	.wren_a(wren_a_1),
	.data_a({a_ram_data_in_bus_59,a_ram_data_in_bus_58,a_ram_data_in_bus_57,a_ram_data_in_bus_56,a_ram_data_in_bus_55,a_ram_data_in_bus_54,a_ram_data_in_bus_53,a_ram_data_in_bus_52,a_ram_data_in_bus_51,a_ram_data_in_bus_50,a_ram_data_in_bus_49,a_ram_data_in_bus_48,
a_ram_data_in_bus_47,a_ram_data_in_bus_46,a_ram_data_in_bus_45,a_ram_data_in_bus_44,a_ram_data_in_bus_43,a_ram_data_in_bus_42,a_ram_data_in_bus_41,a_ram_data_in_bus_40}),
	.clock0(clk));

endmodule

module fftsign_altsyncram_8 (
	q_b,
	clocken0,
	address_a,
	address_b,
	wren_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	wren_a;
input 	[19:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_d0q3_1 auto_generated(
	.q_b({q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clocken0(clocken0),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_d0q3_1 (
	q_b,
	clocken0,
	address_a,
	address_b,
	wren_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	wren_a;
input 	[19:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 20;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 20;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 20;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 20;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 20;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 20;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 20;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 20;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 20;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 20;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 20;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 20;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 20;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "clear0";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "clear0";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 20;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 20;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 20;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 20;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "clear0";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "clear0";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 20;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 20;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 20;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 20;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "clear0";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "clear0";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 20;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 20;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 20;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 20;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "clear0";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "clear0";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 20;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 20;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 20;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 20;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 20;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 20;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 20;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 20;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 20;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 20;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 20;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 20;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 20;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 20;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 20;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module fftsign_asj_fft_data_ram_2 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	wraddress_a_bus_24,
	wraddress_a_bus_10,
	wraddress_a_bus_12,
	rdaddress_a_bus_24,
	rdaddress_a_bus_10,
	rdaddress_a_bus_12,
	rdaddress_a_bus_14,
	wren_a_2,
	a_ram_data_in_bus_32,
	wraddress_a_bus_9,
	wraddress_a_bus_11,
	wraddress_a_bus_13,
	rdaddress_a_bus_9,
	rdaddress_a_bus_11,
	rdaddress_a_bus_13,
	rdaddress_a_bus_15,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_23,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_14;
input 	wren_a_2;
input 	a_ram_data_in_bus_32;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_13;
input 	rdaddress_a_bus_15;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_23;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_dual_port_ram_2 \gen_M4K:ram_component (
	.q_b_12(q_b_12),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_1(q_b_1),
	.q_b_10(q_b_10),
	.q_b_0(q_b_0),
	.q_b_19(q_b_19),
	.q_b_9(q_b_9),
	.q_b_18(q_b_18),
	.q_b_8(q_b_8),
	.q_b_17(q_b_17),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_3(q_b_3),
	.global_clock_enable(global_clock_enable),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.wraddress_a_bus_24(wraddress_a_bus_24),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.rdaddress_a_bus_24(rdaddress_a_bus_24),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_14(rdaddress_a_bus_14),
	.wren_a_2(wren_a_2),
	.a_ram_data_in_bus_32(a_ram_data_in_bus_32),
	.wraddress_a_bus_9(wraddress_a_bus_9),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_9(rdaddress_a_bus_9),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.rdaddress_a_bus_15(rdaddress_a_bus_15),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_39(a_ram_data_in_bus_39),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_38(a_ram_data_in_bus_38),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_37(a_ram_data_in_bus_37),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_36(a_ram_data_in_bus_36),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.a_ram_data_in_bus_35(a_ram_data_in_bus_35),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_34(a_ram_data_in_bus_34),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_33(a_ram_data_in_bus_33),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.clk(clk));

endmodule

module fftsign_altera_fft_dual_port_ram_2 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	wraddress_a_bus_24,
	wraddress_a_bus_10,
	wraddress_a_bus_12,
	rdaddress_a_bus_24,
	rdaddress_a_bus_10,
	rdaddress_a_bus_12,
	rdaddress_a_bus_14,
	wren_a_2,
	a_ram_data_in_bus_32,
	wraddress_a_bus_9,
	wraddress_a_bus_11,
	wraddress_a_bus_13,
	rdaddress_a_bus_9,
	rdaddress_a_bus_11,
	rdaddress_a_bus_13,
	rdaddress_a_bus_15,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_23,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	wraddress_a_bus_24;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_24;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_14;
input 	wren_a_2;
input 	a_ram_data_in_bus_32;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_11;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_11;
input 	rdaddress_a_bus_13;
input 	rdaddress_a_bus_15;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_30;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_23;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_9 \old_ram_gen:old_ram_component (
	.q_b({q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clocken0(global_clock_enable),
	.address_a({wraddress_a_bus_15,wraddress_a_bus_14,wraddress_a_bus_13,wraddress_a_bus_12,wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_9,wraddress_a_bus_24}),
	.address_b({rdaddress_a_bus_15,rdaddress_a_bus_14,rdaddress_a_bus_13,rdaddress_a_bus_12,rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_9,rdaddress_a_bus_24}),
	.wren_a(wren_a_2),
	.data_a({a_ram_data_in_bus_39,a_ram_data_in_bus_38,a_ram_data_in_bus_37,a_ram_data_in_bus_36,a_ram_data_in_bus_35,a_ram_data_in_bus_34,a_ram_data_in_bus_33,a_ram_data_in_bus_32,a_ram_data_in_bus_31,a_ram_data_in_bus_30,a_ram_data_in_bus_29,a_ram_data_in_bus_28,
a_ram_data_in_bus_27,a_ram_data_in_bus_26,a_ram_data_in_bus_25,a_ram_data_in_bus_24,a_ram_data_in_bus_23,a_ram_data_in_bus_22,a_ram_data_in_bus_21,a_ram_data_in_bus_20}),
	.clock0(clk));

endmodule

module fftsign_altsyncram_9 (
	q_b,
	clocken0,
	address_a,
	address_b,
	wren_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	wren_a;
input 	[19:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_d0q3_2 auto_generated(
	.q_b({q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clocken0(clocken0),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_d0q3_2 (
	q_b,
	clocken0,
	address_a,
	address_b,
	wren_a,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	wren_a;
input 	[19:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 20;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 20;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 20;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 20;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 20;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 20;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 20;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 20;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 20;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 20;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 20;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 20;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 20;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "clear0";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "clear0";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 20;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 20;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 20;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 20;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "clear0";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "clear0";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 20;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 20;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 20;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 20;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "clear0";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "clear0";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 20;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 20;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 20;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 20;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "clear0";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "clear0";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 20;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 20;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 20;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 20;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 20;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 20;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 20;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 20;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 20;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 20;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 20;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 20;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 20;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 20;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 20;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module fftsign_asj_fft_data_ram_3 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wren_a_3,
	a_ram_data_in_bus_12,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_18,
	wraddress_a_bus_3,
	wraddress_a_bus_20,
	wraddress_a_bus_5,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_18,
	rdaddress_a_bus_3,
	rdaddress_a_bus_20,
	rdaddress_a_bus_5,
	rdaddress_a_bus_22,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_3,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wren_a_3;
input 	a_ram_data_in_bus_12;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_20;
input 	wraddress_a_bus_5;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_20;
input 	rdaddress_a_bus_5;
input 	rdaddress_a_bus_22;
input 	rdaddress_a_bus_7;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_dual_port_ram_3 \gen_M4K:ram_component (
	.q_b_12(q_b_12),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_1(q_b_1),
	.q_b_10(q_b_10),
	.q_b_0(q_b_0),
	.q_b_19(q_b_19),
	.q_b_9(q_b_9),
	.q_b_18(q_b_18),
	.q_b_8(q_b_8),
	.q_b_17(q_b_17),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_3(q_b_3),
	.global_clock_enable(global_clock_enable),
	.wren_a_3(wren_a_3),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.wraddress_a_bus_18(wraddress_a_bus_18),
	.wraddress_a_bus_3(wraddress_a_bus_3),
	.wraddress_a_bus_20(wraddress_a_bus_20),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.wraddress_a_bus_14(wraddress_a_bus_14),
	.wraddress_a_bus_15(wraddress_a_bus_15),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.rdaddress_a_bus_18(rdaddress_a_bus_18),
	.rdaddress_a_bus_3(rdaddress_a_bus_3),
	.rdaddress_a_bus_20(rdaddress_a_bus_20),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.rdaddress_a_bus_22(rdaddress_a_bus_22),
	.rdaddress_a_bus_7(rdaddress_a_bus_7),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.clk(clk));

endmodule

module fftsign_altera_fft_dual_port_ram_3 (
	q_b_12,
	q_b_2,
	q_b_11,
	q_b_1,
	q_b_10,
	q_b_0,
	q_b_19,
	q_b_9,
	q_b_18,
	q_b_8,
	q_b_17,
	q_b_7,
	q_b_16,
	q_b_6,
	q_b_15,
	q_b_5,
	q_b_14,
	q_b_4,
	q_b_13,
	q_b_3,
	global_clock_enable,
	wren_a_3,
	a_ram_data_in_bus_12,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_18,
	wraddress_a_bus_3,
	wraddress_a_bus_20,
	wraddress_a_bus_5,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_18,
	rdaddress_a_bus_3,
	rdaddress_a_bus_20,
	rdaddress_a_bus_5,
	rdaddress_a_bus_22,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_3,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_2;
output 	q_b_11;
output 	q_b_1;
output 	q_b_10;
output 	q_b_0;
output 	q_b_19;
output 	q_b_9;
output 	q_b_18;
output 	q_b_8;
output 	q_b_17;
output 	q_b_7;
output 	q_b_16;
output 	q_b_6;
output 	q_b_15;
output 	q_b_5;
output 	q_b_14;
output 	q_b_4;
output 	q_b_13;
output 	q_b_3;
input 	global_clock_enable;
input 	wren_a_3;
input 	a_ram_data_in_bus_12;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_1;
input 	wraddress_a_bus_18;
input 	wraddress_a_bus_3;
input 	wraddress_a_bus_20;
input 	wraddress_a_bus_5;
input 	wraddress_a_bus_14;
input 	wraddress_a_bus_15;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_1;
input 	rdaddress_a_bus_18;
input 	rdaddress_a_bus_3;
input 	rdaddress_a_bus_20;
input 	rdaddress_a_bus_5;
input 	rdaddress_a_bus_22;
input 	rdaddress_a_bus_7;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_17;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_14;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_10 \old_ram_gen:old_ram_component (
	.q_b({q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clocken0(global_clock_enable),
	.wren_a(wren_a_3),
	.data_a({a_ram_data_in_bus_19,a_ram_data_in_bus_18,a_ram_data_in_bus_17,a_ram_data_in_bus_16,a_ram_data_in_bus_15,a_ram_data_in_bus_14,a_ram_data_in_bus_13,a_ram_data_in_bus_12,a_ram_data_in_bus_11,a_ram_data_in_bus_10,a_ram_data_in_bus_9,a_ram_data_in_bus_8,
a_ram_data_in_bus_7,a_ram_data_in_bus_6,a_ram_data_in_bus_5,a_ram_data_in_bus_4,a_ram_data_in_bus_3,a_ram_data_in_bus_2,a_ram_data_in_bus_1,a_ram_data_in_bus_0}),
	.address_a({wraddress_a_bus_15,wraddress_a_bus_14,wraddress_a_bus_5,wraddress_a_bus_20,wraddress_a_bus_3,wraddress_a_bus_18,wraddress_a_bus_1,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_7,rdaddress_a_bus_22,rdaddress_a_bus_5,rdaddress_a_bus_20,rdaddress_a_bus_3,rdaddress_a_bus_18,rdaddress_a_bus_1,rdaddress_a_bus_0}),
	.clock0(clk));

endmodule

module fftsign_altsyncram_10 (
	q_b,
	clocken0,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	wren_a;
input 	[19:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altsyncram_d0q3_3 auto_generated(
	.q_b({q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module fftsign_altsyncram_d0q3_3 (
	q_b,
	clocken0,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	clocken0;
input 	wren_a;
input 	[19:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 20;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 20;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 20;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 20;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 20;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 20;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 20;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 20;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 20;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 20;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 20;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 20;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 20;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "clear0";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "clear0";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 20;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 20;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 20;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 20;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "clear0";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "clear0";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 20;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 20;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 20;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 20;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "clear0";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "clear0";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 20;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 20;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 20;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 20;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "clear0";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "clear0";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 20;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 20;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 20;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 20;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 20;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 20;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 20;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 20;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 20;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 20;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 20;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 20;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 20;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_d0q3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 20;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 20;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module fftsign_asj_fft_bfp_ctrl (
	global_clock_enable,
	stall_reg,
	source_stall_int_d,
	global_clock_enable1,
	blk_exp_0,
	blk_exp_1,
	blk_exp_2,
	blk_exp_3,
	blk_exp_4,
	blk_exp_5,
	exp_en,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	tdl_arr_23,
	Mux1,
	tdl_arr_6,
	tdl_arr_9,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable1;
output 	blk_exp_0;
output 	blk_exp_1;
output 	blk_exp_2;
output 	blk_exp_3;
output 	blk_exp_4;
output 	blk_exp_5;
input 	exp_en;
output 	slb_last_0;
output 	slb_last_1;
output 	slb_last_2;
input 	slb_i_0;
input 	slb_i_1;
input 	slb_i_2;
input 	slb_i_3;
input 	Mux2;
input 	tdl_arr_23;
input 	Mux1;
output 	tdl_arr_6;
input 	tdl_arr_9;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ;
wire \blk_exp_acc[0]~6_combout ;
wire \blk_exp_acc[3]~8_combout ;
wire \blk_exp_acc[0]~9_combout ;
wire \blk_exp_acc[0]~10_combout ;
wire \blk_exp_acc[0]~q ;
wire \blk_exp~0_combout ;
wire \blk_exp[0]~1_combout ;
wire \blk_exp_acc[0]~7 ;
wire \blk_exp_acc[1]~11_combout ;
wire \blk_exp_acc[1]~q ;
wire \blk_exp~2_combout ;
wire \blk_exp_acc[1]~12 ;
wire \blk_exp_acc[2]~13_combout ;
wire \blk_exp_acc[2]~q ;
wire \blk_exp~3_combout ;
wire \blk_exp_acc[2]~14 ;
wire \blk_exp_acc[3]~15_combout ;
wire \blk_exp_acc[3]~q ;
wire \blk_exp~4_combout ;
wire \blk_exp_acc[3]~16 ;
wire \blk_exp_acc[4]~17_combout ;
wire \blk_exp_acc[4]~q ;
wire \blk_exp~5_combout ;
wire \blk_exp_acc[4]~18 ;
wire \blk_exp_acc[5]~19_combout ;
wire \blk_exp_acc[5]~q ;
wire \blk_exp~6_combout ;
wire \slb_last~8_combout ;
wire \slb_last[2]~4_combout ;
wire \slb_last[2]~5_combout ;
wire \slb_last~9_combout ;
wire \slb_last~6_combout ;
wire \slb_last~7_combout ;


fftsign_asj_fft_tdl_bit_rst \gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass (
	.global_clock_enable(global_clock_enable1),
	.tdl_arr_9(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.tdl_arr_6(tdl_arr_6),
	.tdl_arr_91(tdl_arr_9),
	.clk(clk),
	.reset_n(reset_n));

dffeas \blk_exp[0] (
	.clk(clk),
	.d(\blk_exp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_0),
	.prn(vcc));
defparam \blk_exp[0] .is_wysiwyg = "true";
defparam \blk_exp[0] .power_up = "low";

dffeas \blk_exp[1] (
	.clk(clk),
	.d(\blk_exp~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_1),
	.prn(vcc));
defparam \blk_exp[1] .is_wysiwyg = "true";
defparam \blk_exp[1] .power_up = "low";

dffeas \blk_exp[2] (
	.clk(clk),
	.d(\blk_exp~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_2),
	.prn(vcc));
defparam \blk_exp[2] .is_wysiwyg = "true";
defparam \blk_exp[2] .power_up = "low";

dffeas \blk_exp[3] (
	.clk(clk),
	.d(\blk_exp~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_3),
	.prn(vcc));
defparam \blk_exp[3] .is_wysiwyg = "true";
defparam \blk_exp[3] .power_up = "low";

dffeas \blk_exp[4] (
	.clk(clk),
	.d(\blk_exp~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_4),
	.prn(vcc));
defparam \blk_exp[4] .is_wysiwyg = "true";
defparam \blk_exp[4] .power_up = "low";

dffeas \blk_exp[5] (
	.clk(clk),
	.d(\blk_exp~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_5),
	.prn(vcc));
defparam \blk_exp[5] .is_wysiwyg = "true";
defparam \blk_exp[5] .power_up = "low";

dffeas \slb_last[0] (
	.clk(clk),
	.d(\slb_last~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_0),
	.prn(vcc));
defparam \slb_last[0] .is_wysiwyg = "true";
defparam \slb_last[0] .power_up = "low";

dffeas \slb_last[1] (
	.clk(clk),
	.d(\slb_last~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_1),
	.prn(vcc));
defparam \slb_last[1] .is_wysiwyg = "true";
defparam \slb_last[1] .power_up = "low";

dffeas \slb_last[2] (
	.clk(clk),
	.d(\slb_last~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~5_combout ),
	.q(slb_last_2),
	.prn(vcc));
defparam \slb_last[2] .is_wysiwyg = "true";
defparam \slb_last[2] .power_up = "low";

cycloneive_lcell_comb \blk_exp_acc[0]~6 (
	.dataa(\blk_exp_acc[0]~q ),
	.datab(slb_last_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~6_combout ),
	.cout(\blk_exp_acc[0]~7 ));
defparam \blk_exp_acc[0]~6 .lut_mask = 16'h66EE;
defparam \blk_exp_acc[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[3]~8 (
	.dataa(reset_n),
	.datab(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[3]~8_combout ),
	.cout());
defparam \blk_exp_acc[3]~8 .lut_mask = 16'h7777;
defparam \blk_exp_acc[3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[0]~9 (
	.dataa(exp_en),
	.datab(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datac(reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~9_combout ),
	.cout());
defparam \blk_exp_acc[0]~9 .lut_mask = 16'hEFEF;
defparam \blk_exp_acc[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[0]~10 (
	.dataa(source_stall_int_d),
	.datab(global_clock_enable),
	.datac(stall_reg),
	.datad(\blk_exp_acc[0]~9_combout ),
	.cin(gnd),
	.combout(\blk_exp_acc[0]~10_combout ),
	.cout());
defparam \blk_exp_acc[0]~10 .lut_mask = 16'hF7D5;
defparam \blk_exp_acc[0]~10 .sum_lutc_input = "datac";

dffeas \blk_exp_acc[0] (
	.clk(clk),
	.d(\blk_exp_acc[0]~6_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[0]~q ),
	.prn(vcc));
defparam \blk_exp_acc[0] .is_wysiwyg = "true";
defparam \blk_exp_acc[0] .power_up = "low";

cycloneive_lcell_comb \blk_exp~0 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~0_combout ),
	.cout());
defparam \blk_exp~0 .lut_mask = 16'hEEEE;
defparam \blk_exp~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp[0]~1 (
	.dataa(global_clock_enable1),
	.datab(reset_n),
	.datac(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datad(exp_en),
	.cin(gnd),
	.combout(\blk_exp[0]~1_combout ),
	.cout());
defparam \blk_exp[0]~1 .lut_mask = 16'hFFBF;
defparam \blk_exp[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[1]~11 (
	.dataa(\blk_exp_acc[1]~q ),
	.datab(slb_last_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[0]~7 ),
	.combout(\blk_exp_acc[1]~11_combout ),
	.cout(\blk_exp_acc[1]~12 ));
defparam \blk_exp_acc[1]~11 .lut_mask = 16'h967F;
defparam \blk_exp_acc[1]~11 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[1] (
	.clk(clk),
	.d(\blk_exp_acc[1]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[1]~q ),
	.prn(vcc));
defparam \blk_exp_acc[1] .is_wysiwyg = "true";
defparam \blk_exp_acc[1] .power_up = "low";

cycloneive_lcell_comb \blk_exp~2 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~2_combout ),
	.cout());
defparam \blk_exp~2 .lut_mask = 16'hEEEE;
defparam \blk_exp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[2]~13 (
	.dataa(\blk_exp_acc[2]~q ),
	.datab(slb_last_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[1]~12 ),
	.combout(\blk_exp_acc[2]~13_combout ),
	.cout(\blk_exp_acc[2]~14 ));
defparam \blk_exp_acc[2]~13 .lut_mask = 16'h96EF;
defparam \blk_exp_acc[2]~13 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[2] (
	.clk(clk),
	.d(\blk_exp_acc[2]~13_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[2]~q ),
	.prn(vcc));
defparam \blk_exp_acc[2] .is_wysiwyg = "true";
defparam \blk_exp_acc[2] .power_up = "low";

cycloneive_lcell_comb \blk_exp~3 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~3_combout ),
	.cout());
defparam \blk_exp~3 .lut_mask = 16'hEEEE;
defparam \blk_exp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[3]~15 (
	.dataa(\blk_exp_acc[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[2]~14 ),
	.combout(\blk_exp_acc[3]~15_combout ),
	.cout(\blk_exp_acc[3]~16 ));
defparam \blk_exp_acc[3]~15 .lut_mask = 16'h5A5F;
defparam \blk_exp_acc[3]~15 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[3] (
	.clk(clk),
	.d(\blk_exp_acc[3]~15_combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[3]~q ),
	.prn(vcc));
defparam \blk_exp_acc[3] .is_wysiwyg = "true";
defparam \blk_exp_acc[3] .power_up = "low";

cycloneive_lcell_comb \blk_exp~4 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~4_combout ),
	.cout());
defparam \blk_exp~4 .lut_mask = 16'hEEEE;
defparam \blk_exp~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[4]~17 (
	.dataa(\blk_exp_acc[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\blk_exp_acc[3]~16 ),
	.combout(\blk_exp_acc[4]~17_combout ),
	.cout(\blk_exp_acc[4]~18 ));
defparam \blk_exp_acc[4]~17 .lut_mask = 16'h5AAF;
defparam \blk_exp_acc[4]~17 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[4] (
	.clk(clk),
	.d(\blk_exp_acc[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[4]~q ),
	.prn(vcc));
defparam \blk_exp_acc[4] .is_wysiwyg = "true";
defparam \blk_exp_acc[4] .power_up = "low";

cycloneive_lcell_comb \blk_exp~5 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~5_combout ),
	.cout());
defparam \blk_exp~5 .lut_mask = 16'hEEEE;
defparam \blk_exp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \blk_exp_acc[5]~19 (
	.dataa(\blk_exp_acc[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\blk_exp_acc[4]~18 ),
	.combout(\blk_exp_acc[5]~19_combout ),
	.cout());
defparam \blk_exp_acc[5]~19 .lut_mask = 16'h5A5A;
defparam \blk_exp_acc[5]~19 .sum_lutc_input = "cin";

dffeas \blk_exp_acc[5] (
	.clk(clk),
	.d(\blk_exp_acc[5]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[3]~8_combout ),
	.ena(\blk_exp_acc[0]~10_combout ),
	.q(\blk_exp_acc[5]~q ),
	.prn(vcc));
defparam \blk_exp_acc[5] .is_wysiwyg = "true";
defparam \blk_exp_acc[5] .power_up = "low";

cycloneive_lcell_comb \blk_exp~6 (
	.dataa(reset_n),
	.datab(\blk_exp_acc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\blk_exp~6_combout ),
	.cout());
defparam \blk_exp~6 .lut_mask = 16'hEEEE;
defparam \blk_exp~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~8 (
	.dataa(reset_n),
	.datab(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datac(Mux2),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last~8_combout ),
	.cout());
defparam \slb_last~8 .lut_mask = 16'hFEFE;
defparam \slb_last~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last[2]~4 (
	.dataa(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datab(tdl_arr_23),
	.datac(reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last[2]~4_combout ),
	.cout());
defparam \slb_last[2]~4 .lut_mask = 16'hEFEF;
defparam \slb_last[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last[2]~5 (
	.dataa(source_stall_int_d),
	.datab(global_clock_enable),
	.datac(stall_reg),
	.datad(\slb_last[2]~4_combout ),
	.cin(gnd),
	.combout(\slb_last[2]~5_combout ),
	.cout());
defparam \slb_last[2]~5 .lut_mask = 16'hF7D5;
defparam \slb_last[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~9 (
	.dataa(reset_n),
	.datab(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datac(Mux1),
	.datad(gnd),
	.cin(gnd),
	.combout(\slb_last~9_combout ),
	.cout());
defparam \slb_last~9 .lut_mask = 16'hFEFE;
defparam \slb_last~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~6 (
	.dataa(reset_n),
	.datab(\gen_quad_burst_ctrl:gen_se_bfp:gen_4bit_accum:delay_next_pass|tdl_arr[9]~q ),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(\slb_last~6_combout ),
	.cout());
defparam \slb_last~6 .lut_mask = 16'hEFFF;
defparam \slb_last~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_last~7 (
	.dataa(\slb_last~6_combout ),
	.datab(gnd),
	.datac(slb_i_0),
	.datad(slb_i_1),
	.cin(gnd),
	.combout(\slb_last~7_combout ),
	.cout());
defparam \slb_last~7 .lut_mask = 16'hAFFF;
defparam \slb_last~7 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_rst (
	global_clock_enable,
	tdl_arr_9,
	tdl_arr_6,
	tdl_arr_91,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_9;
output 	tdl_arr_6;
input 	tdl_arr_91;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~2_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~0_combout ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~3_combout ;


dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(tdl_arr_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(tdl_arr_91),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_addr (
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_5_0,
	ram_in_reg_6_1,
	ram_in_reg_7_3,
	ram_in_reg_7_2,
	rd_addr_d_0,
	rd_addr_d_1,
	rd_addr_d_2,
	rd_addr_d_3,
	rd_addr_d_4,
	rd_addr_d_5,
	sw_0,
	sw_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_6_1;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_2;
input 	rd_addr_d_0;
input 	rd_addr_d_1;
input 	rd_addr_d_2;
input 	rd_addr_d_3;
input 	rd_addr_d_4;
input 	rd_addr_d_5;
input 	sw_0;
input 	sw_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[1][6]~0_combout ;
wire \ram_in_reg[3][7]~1_combout ;
wire \Mux16~0_combout ;


dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(rd_addr_d_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(rd_addr_d_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(rd_addr_d_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(rd_addr_d_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(rd_addr_d_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(rd_addr_d_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\Mux16~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

cycloneive_lcell_comb \ram_in_reg[1][6]~0 (
	.dataa(sw_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~0_combout ),
	.cout());
defparam \ram_in_reg[1][6]~0 .lut_mask = 16'h5555;
defparam \ram_in_reg[1][6]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][7]~1 (
	.dataa(sw_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~1_combout ),
	.cout());
defparam \ram_in_reg[3][7]~1 .lut_mask = 16'h5555;
defparam \ram_in_reg[3][7]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'h0FF0;
defparam \Mux16~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_addr_1 (
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_1,
	ram_in_reg_3_3,
	ram_in_reg_4_1,
	ram_in_reg_5_3,
	ram_in_reg_6_0,
	ram_in_reg_7_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_5_0,
	ram_in_reg_1_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_1_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	rd_addr_c_0,
	rd_addr_d_0,
	sw_0,
	rd_addr_b_1,
	rd_addr_d_1,
	sw_1,
	rd_addr_c_2,
	rd_addr_d_2,
	rd_addr_b_3,
	rd_addr_d_3,
	rd_addr_c_4,
	rd_addr_d_4,
	rd_addr_b_5,
	rd_addr_d_5,
	rd_addr_d_6,
	rd_addr_d_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_3;
output 	ram_in_reg_2_1;
output 	ram_in_reg_3_3;
output 	ram_in_reg_4_1;
output 	ram_in_reg_5_3;
output 	ram_in_reg_6_0;
output 	ram_in_reg_7_0;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_1_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_5_2;
input 	rd_addr_c_0;
input 	rd_addr_d_0;
input 	sw_0;
input 	rd_addr_b_1;
input 	rd_addr_d_1;
input 	sw_1;
input 	rd_addr_c_2;
input 	rd_addr_d_2;
input 	rd_addr_b_3;
input 	rd_addr_d_3;
input 	rd_addr_c_4;
input 	rd_addr_d_4;
input 	rd_addr_b_5;
input 	rd_addr_d_5;
input 	rd_addr_d_6;
input 	rd_addr_d_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux15~0_combout ;
wire \Mux6~0_combout ;
wire \Mux13~0_combout ;
wire \Mux4~0_combout ;
wire \Mux11~0_combout ;
wire \Mux2~0_combout ;
wire \Mux7~0_combout ;
wire \Mux6~1_combout ;
wire \Mux5~0_combout ;
wire \Mux4~1_combout ;
wire \Mux3~0_combout ;
wire \Mux2~1_combout ;
wire \Mux6~2_combout ;
wire \Mux4~2_combout ;
wire \Mux2~2_combout ;
wire \Mux22~0_combout ;
wire \Mux20~0_combout ;
wire \Mux18~0_combout ;


dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(rd_addr_d_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(rd_addr_d_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux4~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux22~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux20~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(rd_addr_c_0),
	.datab(rd_addr_d_0),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAACC;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(rd_addr_b_1),
	.datab(rd_addr_d_1),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hAACC;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(rd_addr_c_2),
	.datab(rd_addr_d_2),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hAACC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(rd_addr_b_3),
	.datab(rd_addr_d_3),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hAACC;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(rd_addr_c_4),
	.datab(rd_addr_d_4),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAACC;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(rd_addr_b_5),
	.datab(rd_addr_d_5),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hAACC;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(rd_addr_d_0),
	.datab(rd_addr_c_0),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hAACC;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(rd_addr_b_1),
	.datab(rd_addr_d_1),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hEFFE;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(rd_addr_d_2),
	.datab(rd_addr_c_2),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hAACC;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(rd_addr_b_3),
	.datab(rd_addr_d_3),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hEFFE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(rd_addr_d_4),
	.datab(rd_addr_c_4),
	.datac(gnd),
	.datad(sw_0),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hAACC;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(rd_addr_b_5),
	.datab(rd_addr_d_5),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hEFFE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(rd_addr_d_1),
	.datab(rd_addr_b_1),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hAACC;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~2 (
	.dataa(rd_addr_d_3),
	.datab(rd_addr_b_3),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
defparam \Mux4~2 .lut_mask = 16'hAACC;
defparam \Mux4~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(rd_addr_d_5),
	.datab(rd_addr_b_5),
	.datac(gnd),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hAACC;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux22~0 (
	.dataa(rd_addr_d_1),
	.datab(rd_addr_b_1),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
defparam \Mux22~0 .lut_mask = 16'hEFFE;
defparam \Mux22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~0 (
	.dataa(rd_addr_d_3),
	.datab(rd_addr_b_3),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
defparam \Mux20~0 .lut_mask = 16'hEFFE;
defparam \Mux20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux18~0 (
	.dataa(rd_addr_d_5),
	.datab(rd_addr_b_5),
	.datac(sw_0),
	.datad(sw_1),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
defparam \Mux18~0 .lut_mask = 16'hEFFE;
defparam \Mux18~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_addr_2 (
	ram_in_reg_1_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	ram_block3a0,
	ram_block3a1,
	ram_in_reg_1_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_1_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_1_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_4_1,
	ram_in_reg_0_11,
	ram_in_reg_1_31,
	ram_in_reg_2_11,
	ram_in_reg_3_31,
	ram_in_reg_4_11,
	ram_in_reg_5_31,
	ram_in_reg_6_0,
	ram_in_reg_7_0,
	ram_in_reg_0_0,
	ram_in_reg_2_0,
	ram_in_reg_4_0,
	ram_in_reg_0_01,
	ram_in_reg_1_01,
	ram_in_reg_2_01,
	ram_in_reg_3_01,
	ram_in_reg_4_01,
	ram_in_reg_5_01,
	ram_in_reg_1_11,
	ram_in_reg_3_11,
	ram_in_reg_5_11,
	ram_in_reg_1_21,
	ram_in_reg_3_21,
	ram_in_reg_5_21,
	swa_tdl_0_16,
	swa_tdl_1_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_1_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_5_3;
output 	ram_block3a0;
output 	ram_block3a1;
output 	ram_in_reg_1_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_1_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_5_2;
input 	global_clock_enable;
output 	ram_in_reg_0_1;
output 	ram_in_reg_2_1;
output 	ram_in_reg_4_1;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_31;
input 	ram_in_reg_2_11;
input 	ram_in_reg_3_31;
input 	ram_in_reg_4_11;
input 	ram_in_reg_5_31;
input 	ram_in_reg_6_0;
input 	ram_in_reg_7_0;
output 	ram_in_reg_0_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_4_0;
input 	ram_in_reg_0_01;
input 	ram_in_reg_1_01;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_4_01;
input 	ram_in_reg_5_01;
input 	ram_in_reg_1_11;
input 	ram_in_reg_3_11;
input 	ram_in_reg_5_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_3_21;
input 	ram_in_reg_5_21;
input 	swa_tdl_0_16;
input 	swa_tdl_1_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ;
wire \ram_in_reg[3][1]~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ;
wire \ram_in_reg[1][1]~6_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10~portbdataout ;
wire \ram_in_reg[3][3]~1_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8~portbdataout ;
wire \ram_in_reg[1][3]~7_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16~portbdataout ;
wire \ram_in_reg[3][5]~2_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14~portbdataout ;
wire \ram_in_reg[1][5]~8_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \ram_in_reg[0][1]~3_combout ;
wire \ram_in_reg[2][1]~9_combout ;
wire \ram_in_reg[0][3]~4_combout ;
wire \ram_in_reg[2][3]~10_combout ;
wire \ram_in_reg[0][5]~5_combout ;
wire \ram_in_reg[2][5]~11_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ;
wire \Mux15~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7~portbdataout ;
wire \Mux13~0_combout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12~portbdataout ;
wire \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13~portbdataout ;
wire \Mux11~0_combout ;
wire \Mux7~0_combout ;
wire \Mux5~0_combout ;
wire \Mux3~0_combout ;

wire [143:0] \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14_PORTBDATAOUT_bus ;

assign ram_block3a0 = \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus [0];

assign ram_block3a1 = \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15_PORTBDATAOUT_bus [0];

assign \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14~portbdataout  = \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14_PORTBDATAOUT_bus [0];

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~0_combout ),
	.asdata(\ram_in_reg[1][1]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~1_combout ),
	.asdata(\ram_in_reg[1][3]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~2_combout ),
	.asdata(\ram_in_reg[1][5]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

cycloneive_ram_block \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_6_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_0|shift_taps_pnm:auto_generated|altsyncram_2e81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_bit_number = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_last_address = 14;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_depth = 15;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_bit_number = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_last_address = 14;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_depth = 15;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a0 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_7_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_0|shift_taps_pnm:auto_generated|altsyncram_2e81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_bit_number = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_last_address = 14;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_depth = 15;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_bit_number = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_last_address = 14;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_depth = 15;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram2|ram_block3a1 .ram_block_type = "auto";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~3_combout ),
	.asdata(\ram_in_reg[2][1]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~4_combout ),
	.asdata(\ram_in_reg[2][3]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~5_combout ),
	.asdata(\ram_in_reg[2][5]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~6_combout ),
	.asdata(\ram_in_reg[3][1]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~7_combout ),
	.asdata(\ram_in_reg[3][3]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~8_combout ),
	.asdata(\ram_in_reg[3][5]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~9_combout ),
	.asdata(\ram_in_reg[0][1]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~10_combout ),
	.asdata(\ram_in_reg[0][3]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~11_combout ),
	.asdata(\ram_in_reg[0][5]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(swa_tdl_1_16),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~combout ),
	.cout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~COUT ));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~combout ),
	.cout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~COUT ));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datac(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datad(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 .lut_mask = 16'hFEFF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~combout ),
	.cout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~COUT ));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~combout ),
	.cout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~COUT ));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 16'h5A5F;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0 .lut_mask = 16'h0F0F;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita0~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_1|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_31}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_first_bit_number = 5;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_first_bit_number = 5;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_21}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_first_bit_number = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_first_bit_number = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[3][1]~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~0_combout ),
	.cout());
defparam \ram_in_reg[3][1]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~0 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_first_bit_number = 3;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_first_bit_number = 3;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_first_bit_number = 2;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_first_bit_number = 2;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[1][1]~6 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~6_combout ),
	.cout());
defparam \ram_in_reg[1][1]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~6 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_3_31}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_first_bit_number = 11;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_first_bit_number = 11;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_3_21}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_first_bit_number = 10;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_first_bit_number = 10;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[3][3]~1 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~1_combout ),
	.cout());
defparam \ram_in_reg[3][3]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~1 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_3_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_first_bit_number = 9;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_first_bit_number = 9;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_3_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_first_bit_number = 8;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_first_bit_number = 8;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[1][3]~7 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~7_combout ),
	.cout());
defparam \ram_in_reg[1][3]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~7 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_5_31}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_first_bit_number = 17;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_first_bit_number = 17;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_5_21}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_first_bit_number = 16;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_first_bit_number = 16;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[3][5]~2 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~2_combout ),
	.cout());
defparam \ram_in_reg[3][5]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~2 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_5_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_first_bit_number = 15;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_first_bit_number = 15;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_5_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_first_bit_number = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_first_bit_number = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14 .ram_block_type = "auto";

cycloneive_lcell_comb \ram_in_reg[1][5]~8 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~8_combout ),
	.cout());
defparam \ram_in_reg[1][5]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datac(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datad(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 .lut_mask = 16'hFEFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 16'h5A5F;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0 .lut_mask = 16'h0F0F;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0 .sum_lutc_input = "cin";

cycloneive_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0 (
	.dataa(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ),
	.datab(gnd),
	.datac(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~0_combout ),
	.datad(\sw_0_arr_rtl_0|auto_generated|cntr1|cmpr4|aneb_result_wire[0]~0_combout ),
	.cin(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0_combout ),
	.cout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0 .lut_mask = 16'hAFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0 .sum_lutc_input = "datac";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb \ram_in_reg[0][1]~3 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a2~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a5~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~3_combout ),
	.cout());
defparam \ram_in_reg[0][1]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][1]~9 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a4~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a3~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~9_combout ),
	.cout());
defparam \ram_in_reg[2][1]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][3]~4 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a8~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a11~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~4_combout ),
	.cout());
defparam \ram_in_reg[0][3]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][3]~10 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a10~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a9~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~10_combout ),
	.cout());
defparam \ram_in_reg[2][3]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][5]~5 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a14~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a17~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~5_combout ),
	.cout());
defparam \ram_in_reg[0][5]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][5]~11 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a16~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a15~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~11_combout ),
	.cout());
defparam \ram_in_reg[2][5]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~11 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_0_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_first_bit_number = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_first_bit_number = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_0_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_first_bit_number = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_first_bit_number = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1 .ram_block_type = "auto";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAACC;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_2_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_first_bit_number = 6;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_first_bit_number = 6;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_2_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_first_bit_number = 7;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_first_bit_number = 7;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7 .ram_block_type = "auto";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hAACC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_4_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_first_bit_number = 12;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_first_bit_number = 12;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12 .ram_block_type = "auto";

cycloneive_ram_block \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_4_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_0_arr_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13_PORTBDATAOUT_bus ));
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .clk0_output_clock_enable = "ena0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_cxb_addr:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_1|shift_taps_fpm:auto_generated|altsyncram_eh81:altsyncram2|ALTSYNCRAM";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .mixed_port_feed_through_mode = "old";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_first_bit_number = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_address_width = 4;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_data_out_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_first_bit_number = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_last_address = 13;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_logical_ram_depth = 14;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_logical_ram_width = 18;
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13 .ram_block_type = "auto";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAACC;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a1~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a0~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hAACC;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a7~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a6~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hAACC;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a13~portbdataout ),
	.datab(\sw_0_arr_rtl_1|auto_generated|altsyncram2|ram_block3a12~portbdataout ),
	.datac(gnd),
	.datad(swa_tdl_0_16),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hAACC;
defparam \Mux3~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_data (
	ram_in_reg_2_3,
	ram_in_reg_2_0,
	ram_in_reg_2_1,
	ram_in_reg_2_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_1_3,
	ram_in_reg_1_0,
	ram_in_reg_1_1,
	ram_in_reg_1_2,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	ram_in_reg_0_3,
	ram_in_reg_0_0,
	ram_in_reg_0_1,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	ram_in_reg_9_3,
	ram_in_reg_9_0,
	ram_in_reg_9_1,
	ram_in_reg_9_2,
	ram_in_reg_9_7,
	ram_in_reg_9_4,
	ram_in_reg_9_5,
	ram_in_reg_9_6,
	ram_in_reg_8_3,
	ram_in_reg_8_0,
	ram_in_reg_8_1,
	ram_in_reg_8_2,
	ram_in_reg_8_7,
	ram_in_reg_8_4,
	ram_in_reg_8_5,
	ram_in_reg_8_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_5_3,
	ram_in_reg_5_0,
	ram_in_reg_5_1,
	ram_in_reg_5_2,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	ram_in_reg_3_1,
	ram_in_reg_3_2,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	ram_block3a1,
	ram_block3a0,
	global_clock_enable,
	reg_no_twiddle605,
	reg_no_twiddle609,
	reg_no_twiddle615,
	reg_no_twiddle619,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_5_12,
	tdl_arr_9_12,
	tdl_arr_5_13,
	tdl_arr_9_13,
	tdl_arr_5_14,
	tdl_arr_9_14,
	tdl_arr_5_15,
	tdl_arr_9_15,
	reg_no_twiddle606,
	reg_no_twiddle616,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	reg_no_twiddle607,
	reg_no_twiddle617,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_7_12,
	tdl_arr_7_13,
	tdl_arr_7_14,
	tdl_arr_7_15,
	reg_no_twiddle608,
	reg_no_twiddle618,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_8_12,
	tdl_arr_8_13,
	tdl_arr_8_14,
	tdl_arr_8_15,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_2_12,
	reg_no_twiddle602,
	tdl_arr_2_13,
	tdl_arr_2_14,
	tdl_arr_2_15,
	reg_no_twiddle612,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_1_12,
	reg_no_twiddle601,
	tdl_arr_1_13,
	tdl_arr_1_14,
	tdl_arr_1_15,
	reg_no_twiddle611,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_0_12,
	reg_no_twiddle600,
	tdl_arr_0_13,
	tdl_arr_0_14,
	tdl_arr_0_15,
	reg_no_twiddle610,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_4_12,
	reg_no_twiddle604,
	tdl_arr_4_13,
	tdl_arr_4_14,
	tdl_arr_4_15,
	reg_no_twiddle614,
	tdl_arr_3_1,
	tdl_arr_3_11,
	tdl_arr_3_12,
	reg_no_twiddle603,
	tdl_arr_3_13,
	tdl_arr_3_14,
	tdl_arr_3_15,
	reg_no_twiddle613,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_2_3;
output 	ram_in_reg_2_0;
output 	ram_in_reg_2_1;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_4;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_6;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_7;
output 	ram_in_reg_1_4;
output 	ram_in_reg_1_5;
output 	ram_in_reg_1_6;
output 	ram_in_reg_0_3;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_7;
output 	ram_in_reg_0_4;
output 	ram_in_reg_0_5;
output 	ram_in_reg_0_6;
output 	ram_in_reg_9_3;
output 	ram_in_reg_9_0;
output 	ram_in_reg_9_1;
output 	ram_in_reg_9_2;
output 	ram_in_reg_9_7;
output 	ram_in_reg_9_4;
output 	ram_in_reg_9_5;
output 	ram_in_reg_9_6;
output 	ram_in_reg_8_3;
output 	ram_in_reg_8_0;
output 	ram_in_reg_8_1;
output 	ram_in_reg_8_2;
output 	ram_in_reg_8_7;
output 	ram_in_reg_8_4;
output 	ram_in_reg_8_5;
output 	ram_in_reg_8_6;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_7;
output 	ram_in_reg_7_4;
output 	ram_in_reg_7_5;
output 	ram_in_reg_7_6;
output 	ram_in_reg_6_3;
output 	ram_in_reg_6_0;
output 	ram_in_reg_6_1;
output 	ram_in_reg_6_2;
output 	ram_in_reg_6_7;
output 	ram_in_reg_6_4;
output 	ram_in_reg_6_5;
output 	ram_in_reg_6_6;
output 	ram_in_reg_5_3;
output 	ram_in_reg_5_0;
output 	ram_in_reg_5_1;
output 	ram_in_reg_5_2;
output 	ram_in_reg_5_7;
output 	ram_in_reg_5_4;
output 	ram_in_reg_5_5;
output 	ram_in_reg_5_6;
output 	ram_in_reg_4_3;
output 	ram_in_reg_4_0;
output 	ram_in_reg_4_1;
output 	ram_in_reg_4_2;
output 	ram_in_reg_4_7;
output 	ram_in_reg_4_4;
output 	ram_in_reg_4_5;
output 	ram_in_reg_4_6;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_0;
output 	ram_in_reg_3_1;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_7;
output 	ram_in_reg_3_4;
output 	ram_in_reg_3_5;
output 	ram_in_reg_3_6;
input 	ram_block3a1;
input 	ram_block3a0;
input 	global_clock_enable;
input 	reg_no_twiddle605;
input 	reg_no_twiddle609;
input 	reg_no_twiddle615;
input 	reg_no_twiddle619;
input 	tdl_arr_5_1;
input 	tdl_arr_9_1;
input 	tdl_arr_5_11;
input 	tdl_arr_9_11;
input 	tdl_arr_5_12;
input 	tdl_arr_9_12;
input 	tdl_arr_5_13;
input 	tdl_arr_9_13;
input 	tdl_arr_5_14;
input 	tdl_arr_9_14;
input 	tdl_arr_5_15;
input 	tdl_arr_9_15;
input 	reg_no_twiddle606;
input 	reg_no_twiddle616;
input 	tdl_arr_6_1;
input 	tdl_arr_6_11;
input 	tdl_arr_6_12;
input 	tdl_arr_6_13;
input 	tdl_arr_6_14;
input 	tdl_arr_6_15;
input 	reg_no_twiddle607;
input 	reg_no_twiddle617;
input 	tdl_arr_7_1;
input 	tdl_arr_7_11;
input 	tdl_arr_7_12;
input 	tdl_arr_7_13;
input 	tdl_arr_7_14;
input 	tdl_arr_7_15;
input 	reg_no_twiddle608;
input 	reg_no_twiddle618;
input 	tdl_arr_8_1;
input 	tdl_arr_8_11;
input 	tdl_arr_8_12;
input 	tdl_arr_8_13;
input 	tdl_arr_8_14;
input 	tdl_arr_8_15;
input 	tdl_arr_2_1;
input 	tdl_arr_2_11;
input 	tdl_arr_2_12;
input 	reg_no_twiddle602;
input 	tdl_arr_2_13;
input 	tdl_arr_2_14;
input 	tdl_arr_2_15;
input 	reg_no_twiddle612;
input 	tdl_arr_1_1;
input 	tdl_arr_1_11;
input 	tdl_arr_1_12;
input 	reg_no_twiddle601;
input 	tdl_arr_1_13;
input 	tdl_arr_1_14;
input 	tdl_arr_1_15;
input 	reg_no_twiddle611;
input 	tdl_arr_0_1;
input 	tdl_arr_0_11;
input 	tdl_arr_0_12;
input 	reg_no_twiddle600;
input 	tdl_arr_0_13;
input 	tdl_arr_0_14;
input 	tdl_arr_0_15;
input 	reg_no_twiddle610;
input 	tdl_arr_4_1;
input 	tdl_arr_4_11;
input 	tdl_arr_4_12;
input 	reg_no_twiddle604;
input 	tdl_arr_4_13;
input 	tdl_arr_4_14;
input 	tdl_arr_4_15;
input 	reg_no_twiddle614;
input 	tdl_arr_3_1;
input 	tdl_arr_3_11;
input 	tdl_arr_3_12;
input 	reg_no_twiddle603;
input 	tdl_arr_3_13;
input 	tdl_arr_3_14;
input 	tdl_arr_3_15;
input 	reg_no_twiddle613;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[3][2]~0_combout ;
wire \ram_in_reg[1][2]~2_combout ;
wire \ram_in_reg[0][2]~1_combout ;
wire \ram_in_reg[2][2]~3_combout ;
wire \ram_in_reg[7][2]~4_combout ;
wire \ram_in_reg[5][2]~6_combout ;
wire \ram_in_reg[4][2]~5_combout ;
wire \ram_in_reg[6][2]~7_combout ;
wire \ram_in_reg[3][1]~64_combout ;
wire \ram_in_reg[1][1]~66_combout ;
wire \ram_in_reg[0][1]~65_combout ;
wire \ram_in_reg[2][1]~67_combout ;
wire \ram_in_reg[7][1]~68_combout ;
wire \ram_in_reg[5][1]~70_combout ;
wire \ram_in_reg[4][1]~69_combout ;
wire \ram_in_reg[6][1]~71_combout ;
wire \ram_in_reg[3][0]~72_combout ;
wire \ram_in_reg[1][0]~74_combout ;
wire \ram_in_reg[0][0]~73_combout ;
wire \ram_in_reg[2][0]~75_combout ;
wire \ram_in_reg[7][0]~76_combout ;
wire \ram_in_reg[5][0]~78_combout ;
wire \ram_in_reg[4][0]~77_combout ;
wire \ram_in_reg[6][0]~79_combout ;
wire \ram_in_reg[3][9]~56_combout ;
wire \ram_in_reg[1][9]~58_combout ;
wire \ram_in_reg[0][9]~57_combout ;
wire \ram_in_reg[2][9]~59_combout ;
wire \ram_in_reg[7][9]~60_combout ;
wire \ram_in_reg[5][9]~62_combout ;
wire \ram_in_reg[4][9]~61_combout ;
wire \ram_in_reg[6][9]~63_combout ;
wire \ram_in_reg[3][8]~48_combout ;
wire \ram_in_reg[1][8]~50_combout ;
wire \ram_in_reg[0][8]~49_combout ;
wire \ram_in_reg[2][8]~51_combout ;
wire \ram_in_reg[7][8]~52_combout ;
wire \ram_in_reg[5][8]~54_combout ;
wire \ram_in_reg[4][8]~53_combout ;
wire \ram_in_reg[6][8]~55_combout ;
wire \ram_in_reg[3][7]~40_combout ;
wire \ram_in_reg[1][7]~42_combout ;
wire \ram_in_reg[0][7]~41_combout ;
wire \ram_in_reg[2][7]~43_combout ;
wire \ram_in_reg[7][7]~44_combout ;
wire \ram_in_reg[5][7]~46_combout ;
wire \ram_in_reg[4][7]~45_combout ;
wire \ram_in_reg[6][7]~47_combout ;
wire \ram_in_reg[3][6]~32_combout ;
wire \ram_in_reg[1][6]~34_combout ;
wire \ram_in_reg[0][6]~33_combout ;
wire \ram_in_reg[2][6]~35_combout ;
wire \ram_in_reg[7][6]~36_combout ;
wire \ram_in_reg[5][6]~38_combout ;
wire \ram_in_reg[4][6]~37_combout ;
wire \ram_in_reg[6][6]~39_combout ;
wire \ram_in_reg[3][5]~24_combout ;
wire \ram_in_reg[1][5]~26_combout ;
wire \ram_in_reg[0][5]~25_combout ;
wire \ram_in_reg[2][5]~27_combout ;
wire \ram_in_reg[7][5]~28_combout ;
wire \ram_in_reg[5][5]~30_combout ;
wire \ram_in_reg[4][5]~29_combout ;
wire \ram_in_reg[6][5]~31_combout ;
wire \ram_in_reg[3][4]~16_combout ;
wire \ram_in_reg[1][4]~18_combout ;
wire \ram_in_reg[0][4]~17_combout ;
wire \ram_in_reg[2][4]~19_combout ;
wire \ram_in_reg[7][4]~20_combout ;
wire \ram_in_reg[5][4]~22_combout ;
wire \ram_in_reg[4][4]~21_combout ;
wire \ram_in_reg[6][4]~23_combout ;
wire \ram_in_reg[3][3]~8_combout ;
wire \ram_in_reg[1][3]~10_combout ;
wire \ram_in_reg[0][3]~9_combout ;
wire \ram_in_reg[2][3]~11_combout ;
wire \ram_in_reg[7][3]~12_combout ;
wire \ram_in_reg[5][3]~14_combout ;
wire \ram_in_reg[4][3]~13_combout ;
wire \ram_in_reg[6][3]~15_combout ;


dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\ram_in_reg[3][2]~0_combout ),
	.asdata(\ram_in_reg[1][2]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\ram_in_reg[0][2]~1_combout ),
	.asdata(\ram_in_reg[2][2]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~2_combout ),
	.asdata(\ram_in_reg[3][2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\ram_in_reg[2][2]~3_combout ),
	.asdata(\ram_in_reg[0][2]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\ram_in_reg[7][2]~4_combout ),
	.asdata(\ram_in_reg[5][2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\ram_in_reg[4][2]~5_combout ),
	.asdata(\ram_in_reg[6][2]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\ram_in_reg[5][2]~6_combout ),
	.asdata(\ram_in_reg[7][2]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\ram_in_reg[6][2]~7_combout ),
	.asdata(\ram_in_reg[4][2]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~64_combout ),
	.asdata(\ram_in_reg[1][1]~66_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~65_combout ),
	.asdata(\ram_in_reg[2][1]~67_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~66_combout ),
	.asdata(\ram_in_reg[3][1]~64_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~67_combout ),
	.asdata(\ram_in_reg[0][1]~65_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\ram_in_reg[7][1]~68_combout ),
	.asdata(\ram_in_reg[5][1]~70_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\ram_in_reg[4][1]~69_combout ),
	.asdata(\ram_in_reg[6][1]~71_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\ram_in_reg[5][1]~70_combout ),
	.asdata(\ram_in_reg[7][1]~68_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\ram_in_reg[6][1]~71_combout ),
	.asdata(\ram_in_reg[4][1]~69_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\ram_in_reg[3][0]~72_combout ),
	.asdata(\ram_in_reg[1][0]~74_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\ram_in_reg[0][0]~73_combout ),
	.asdata(\ram_in_reg[2][0]~75_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\ram_in_reg[1][0]~74_combout ),
	.asdata(\ram_in_reg[3][0]~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\ram_in_reg[2][0]~75_combout ),
	.asdata(\ram_in_reg[0][0]~73_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\ram_in_reg[7][0]~76_combout ),
	.asdata(\ram_in_reg[5][0]~78_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\ram_in_reg[4][0]~77_combout ),
	.asdata(\ram_in_reg[6][0]~79_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\ram_in_reg[5][0]~78_combout ),
	.asdata(\ram_in_reg[7][0]~76_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\ram_in_reg[6][0]~79_combout ),
	.asdata(\ram_in_reg[4][0]~77_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[3][9] (
	.clk(clk),
	.d(\ram_in_reg[3][9]~56_combout ),
	.asdata(\ram_in_reg[1][9]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_3),
	.prn(vcc));
defparam \ram_in_reg[3][9] .is_wysiwyg = "true";
defparam \ram_in_reg[3][9] .power_up = "low";

dffeas \ram_in_reg[0][9] (
	.clk(clk),
	.d(\ram_in_reg[0][9]~57_combout ),
	.asdata(\ram_in_reg[2][9]~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_0),
	.prn(vcc));
defparam \ram_in_reg[0][9] .is_wysiwyg = "true";
defparam \ram_in_reg[0][9] .power_up = "low";

dffeas \ram_in_reg[1][9] (
	.clk(clk),
	.d(\ram_in_reg[1][9]~58_combout ),
	.asdata(\ram_in_reg[3][9]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_1),
	.prn(vcc));
defparam \ram_in_reg[1][9] .is_wysiwyg = "true";
defparam \ram_in_reg[1][9] .power_up = "low";

dffeas \ram_in_reg[2][9] (
	.clk(clk),
	.d(\ram_in_reg[2][9]~59_combout ),
	.asdata(\ram_in_reg[0][9]~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_2),
	.prn(vcc));
defparam \ram_in_reg[2][9] .is_wysiwyg = "true";
defparam \ram_in_reg[2][9] .power_up = "low";

dffeas \ram_in_reg[7][9] (
	.clk(clk),
	.d(\ram_in_reg[7][9]~60_combout ),
	.asdata(\ram_in_reg[5][9]~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_7),
	.prn(vcc));
defparam \ram_in_reg[7][9] .is_wysiwyg = "true";
defparam \ram_in_reg[7][9] .power_up = "low";

dffeas \ram_in_reg[4][9] (
	.clk(clk),
	.d(\ram_in_reg[4][9]~61_combout ),
	.asdata(\ram_in_reg[6][9]~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_4),
	.prn(vcc));
defparam \ram_in_reg[4][9] .is_wysiwyg = "true";
defparam \ram_in_reg[4][9] .power_up = "low";

dffeas \ram_in_reg[5][9] (
	.clk(clk),
	.d(\ram_in_reg[5][9]~62_combout ),
	.asdata(\ram_in_reg[7][9]~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_5),
	.prn(vcc));
defparam \ram_in_reg[5][9] .is_wysiwyg = "true";
defparam \ram_in_reg[5][9] .power_up = "low";

dffeas \ram_in_reg[6][9] (
	.clk(clk),
	.d(\ram_in_reg[6][9]~63_combout ),
	.asdata(\ram_in_reg[4][9]~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_6),
	.prn(vcc));
defparam \ram_in_reg[6][9] .is_wysiwyg = "true";
defparam \ram_in_reg[6][9] .power_up = "low";

dffeas \ram_in_reg[3][8] (
	.clk(clk),
	.d(\ram_in_reg[3][8]~48_combout ),
	.asdata(\ram_in_reg[1][8]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_3),
	.prn(vcc));
defparam \ram_in_reg[3][8] .is_wysiwyg = "true";
defparam \ram_in_reg[3][8] .power_up = "low";

dffeas \ram_in_reg[0][8] (
	.clk(clk),
	.d(\ram_in_reg[0][8]~49_combout ),
	.asdata(\ram_in_reg[2][8]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_0),
	.prn(vcc));
defparam \ram_in_reg[0][8] .is_wysiwyg = "true";
defparam \ram_in_reg[0][8] .power_up = "low";

dffeas \ram_in_reg[1][8] (
	.clk(clk),
	.d(\ram_in_reg[1][8]~50_combout ),
	.asdata(\ram_in_reg[3][8]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_1),
	.prn(vcc));
defparam \ram_in_reg[1][8] .is_wysiwyg = "true";
defparam \ram_in_reg[1][8] .power_up = "low";

dffeas \ram_in_reg[2][8] (
	.clk(clk),
	.d(\ram_in_reg[2][8]~51_combout ),
	.asdata(\ram_in_reg[0][8]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_2),
	.prn(vcc));
defparam \ram_in_reg[2][8] .is_wysiwyg = "true";
defparam \ram_in_reg[2][8] .power_up = "low";

dffeas \ram_in_reg[7][8] (
	.clk(clk),
	.d(\ram_in_reg[7][8]~52_combout ),
	.asdata(\ram_in_reg[5][8]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_7),
	.prn(vcc));
defparam \ram_in_reg[7][8] .is_wysiwyg = "true";
defparam \ram_in_reg[7][8] .power_up = "low";

dffeas \ram_in_reg[4][8] (
	.clk(clk),
	.d(\ram_in_reg[4][8]~53_combout ),
	.asdata(\ram_in_reg[6][8]~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_4),
	.prn(vcc));
defparam \ram_in_reg[4][8] .is_wysiwyg = "true";
defparam \ram_in_reg[4][8] .power_up = "low";

dffeas \ram_in_reg[5][8] (
	.clk(clk),
	.d(\ram_in_reg[5][8]~54_combout ),
	.asdata(\ram_in_reg[7][8]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_5),
	.prn(vcc));
defparam \ram_in_reg[5][8] .is_wysiwyg = "true";
defparam \ram_in_reg[5][8] .power_up = "low";

dffeas \ram_in_reg[6][8] (
	.clk(clk),
	.d(\ram_in_reg[6][8]~55_combout ),
	.asdata(\ram_in_reg[4][8]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_6),
	.prn(vcc));
defparam \ram_in_reg[6][8] .is_wysiwyg = "true";
defparam \ram_in_reg[6][8] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~40_combout ),
	.asdata(\ram_in_reg[1][7]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\ram_in_reg[0][7]~41_combout ),
	.asdata(\ram_in_reg[2][7]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\ram_in_reg[1][7]~42_combout ),
	.asdata(\ram_in_reg[3][7]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\ram_in_reg[2][7]~43_combout ),
	.asdata(\ram_in_reg[0][7]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\ram_in_reg[7][7]~44_combout ),
	.asdata(\ram_in_reg[5][7]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\ram_in_reg[4][7]~45_combout ),
	.asdata(\ram_in_reg[6][7]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\ram_in_reg[5][7]~46_combout ),
	.asdata(\ram_in_reg[7][7]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\ram_in_reg[6][7]~47_combout ),
	.asdata(\ram_in_reg[4][7]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\ram_in_reg[3][6]~32_combout ),
	.asdata(\ram_in_reg[1][6]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\ram_in_reg[0][6]~33_combout ),
	.asdata(\ram_in_reg[2][6]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~34_combout ),
	.asdata(\ram_in_reg[3][6]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\ram_in_reg[2][6]~35_combout ),
	.asdata(\ram_in_reg[0][6]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\ram_in_reg[7][6]~36_combout ),
	.asdata(\ram_in_reg[5][6]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\ram_in_reg[4][6]~37_combout ),
	.asdata(\ram_in_reg[6][6]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\ram_in_reg[5][6]~38_combout ),
	.asdata(\ram_in_reg[7][6]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\ram_in_reg[6][6]~39_combout ),
	.asdata(\ram_in_reg[4][6]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~24_combout ),
	.asdata(\ram_in_reg[1][5]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~25_combout ),
	.asdata(\ram_in_reg[2][5]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~26_combout ),
	.asdata(\ram_in_reg[3][5]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~27_combout ),
	.asdata(\ram_in_reg[0][5]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\ram_in_reg[7][5]~28_combout ),
	.asdata(\ram_in_reg[5][5]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\ram_in_reg[4][5]~29_combout ),
	.asdata(\ram_in_reg[6][5]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\ram_in_reg[5][5]~30_combout ),
	.asdata(\ram_in_reg[7][5]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\ram_in_reg[6][5]~31_combout ),
	.asdata(\ram_in_reg[4][5]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\ram_in_reg[3][4]~16_combout ),
	.asdata(\ram_in_reg[1][4]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\ram_in_reg[0][4]~17_combout ),
	.asdata(\ram_in_reg[2][4]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\ram_in_reg[1][4]~18_combout ),
	.asdata(\ram_in_reg[3][4]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\ram_in_reg[2][4]~19_combout ),
	.asdata(\ram_in_reg[0][4]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\ram_in_reg[7][4]~20_combout ),
	.asdata(\ram_in_reg[5][4]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\ram_in_reg[4][4]~21_combout ),
	.asdata(\ram_in_reg[6][4]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\ram_in_reg[5][4]~22_combout ),
	.asdata(\ram_in_reg[7][4]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\ram_in_reg[6][4]~23_combout ),
	.asdata(\ram_in_reg[4][4]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~8_combout ),
	.asdata(\ram_in_reg[1][3]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~9_combout ),
	.asdata(\ram_in_reg[2][3]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~10_combout ),
	.asdata(\ram_in_reg[3][3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~11_combout ),
	.asdata(\ram_in_reg[0][3]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\ram_in_reg[7][3]~12_combout ),
	.asdata(\ram_in_reg[5][3]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\ram_in_reg[4][3]~13_combout ),
	.asdata(\ram_in_reg[6][3]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\ram_in_reg[5][3]~14_combout ),
	.asdata(\ram_in_reg[7][3]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\ram_in_reg[6][3]~15_combout ),
	.asdata(\ram_in_reg[4][3]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(ram_block3a0),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

cycloneive_lcell_comb \ram_in_reg[3][2]~0 (
	.dataa(tdl_arr_2_1),
	.datab(tdl_arr_2_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][2]~0_combout ),
	.cout());
defparam \ram_in_reg[3][2]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][2]~2 (
	.dataa(tdl_arr_2_12),
	.datab(reg_no_twiddle602),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][2]~2_combout ),
	.cout());
defparam \ram_in_reg[1][2]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][2]~1 (
	.dataa(reg_no_twiddle602),
	.datab(tdl_arr_2_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][2]~1_combout ),
	.cout());
defparam \ram_in_reg[0][2]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][2]~3 (
	.dataa(tdl_arr_2_11),
	.datab(tdl_arr_2_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][2]~3_combout ),
	.cout());
defparam \ram_in_reg[2][2]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][2]~4 (
	.dataa(tdl_arr_2_13),
	.datab(tdl_arr_2_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][2]~4_combout ),
	.cout());
defparam \ram_in_reg[7][2]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][2]~6 (
	.dataa(tdl_arr_2_15),
	.datab(reg_no_twiddle612),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][2]~6_combout ),
	.cout());
defparam \ram_in_reg[5][2]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][2]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][2]~5 (
	.dataa(reg_no_twiddle612),
	.datab(tdl_arr_2_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][2]~5_combout ),
	.cout());
defparam \ram_in_reg[4][2]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][2]~7 (
	.dataa(tdl_arr_2_14),
	.datab(tdl_arr_2_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][2]~7_combout ),
	.cout());
defparam \ram_in_reg[6][2]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][2]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][1]~64 (
	.dataa(tdl_arr_1_1),
	.datab(tdl_arr_1_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~64_combout ),
	.cout());
defparam \ram_in_reg[3][1]~64 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][1]~66 (
	.dataa(tdl_arr_1_12),
	.datab(reg_no_twiddle601),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~66_combout ),
	.cout());
defparam \ram_in_reg[1][1]~66 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][1]~65 (
	.dataa(reg_no_twiddle601),
	.datab(tdl_arr_1_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~65_combout ),
	.cout());
defparam \ram_in_reg[0][1]~65 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][1]~67 (
	.dataa(tdl_arr_1_11),
	.datab(tdl_arr_1_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~67_combout ),
	.cout());
defparam \ram_in_reg[2][1]~67 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][1]~68 (
	.dataa(tdl_arr_1_13),
	.datab(tdl_arr_1_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][1]~68_combout ),
	.cout());
defparam \ram_in_reg[7][1]~68 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][1]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][1]~70 (
	.dataa(tdl_arr_1_15),
	.datab(reg_no_twiddle611),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][1]~70_combout ),
	.cout());
defparam \ram_in_reg[5][1]~70 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][1]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][1]~69 (
	.dataa(reg_no_twiddle611),
	.datab(tdl_arr_1_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][1]~69_combout ),
	.cout());
defparam \ram_in_reg[4][1]~69 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][1]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][1]~71 (
	.dataa(tdl_arr_1_14),
	.datab(tdl_arr_1_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][1]~71_combout ),
	.cout());
defparam \ram_in_reg[6][1]~71 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][1]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][0]~72 (
	.dataa(tdl_arr_0_1),
	.datab(tdl_arr_0_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][0]~72_combout ),
	.cout());
defparam \ram_in_reg[3][0]~72 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][0]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][0]~74 (
	.dataa(tdl_arr_0_12),
	.datab(reg_no_twiddle600),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][0]~74_combout ),
	.cout());
defparam \ram_in_reg[1][0]~74 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][0]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][0]~73 (
	.dataa(reg_no_twiddle600),
	.datab(tdl_arr_0_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][0]~73_combout ),
	.cout());
defparam \ram_in_reg[0][0]~73 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][0]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][0]~75 (
	.dataa(tdl_arr_0_11),
	.datab(tdl_arr_0_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][0]~75_combout ),
	.cout());
defparam \ram_in_reg[2][0]~75 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][0]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][0]~76 (
	.dataa(tdl_arr_0_13),
	.datab(tdl_arr_0_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][0]~76_combout ),
	.cout());
defparam \ram_in_reg[7][0]~76 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][0]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][0]~78 (
	.dataa(tdl_arr_0_15),
	.datab(reg_no_twiddle610),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][0]~78_combout ),
	.cout());
defparam \ram_in_reg[5][0]~78 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][0]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][0]~77 (
	.dataa(reg_no_twiddle610),
	.datab(tdl_arr_0_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][0]~77_combout ),
	.cout());
defparam \ram_in_reg[4][0]~77 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][0]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][0]~79 (
	.dataa(tdl_arr_0_14),
	.datab(tdl_arr_0_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][0]~79_combout ),
	.cout());
defparam \ram_in_reg[6][0]~79 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][0]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][9]~56 (
	.dataa(tdl_arr_9_14),
	.datab(tdl_arr_9_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][9]~56_combout ),
	.cout());
defparam \ram_in_reg[3][9]~56 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][9]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][9]~58 (
	.dataa(tdl_arr_9_1),
	.datab(reg_no_twiddle609),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][9]~58_combout ),
	.cout());
defparam \ram_in_reg[1][9]~58 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][9]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][9]~57 (
	.dataa(reg_no_twiddle609),
	.datab(tdl_arr_9_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][9]~57_combout ),
	.cout());
defparam \ram_in_reg[0][9]~57 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][9]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][9]~59 (
	.dataa(tdl_arr_9_12),
	.datab(tdl_arr_9_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][9]~59_combout ),
	.cout());
defparam \ram_in_reg[2][9]~59 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][9]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][9]~60 (
	.dataa(tdl_arr_9_15),
	.datab(tdl_arr_9_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][9]~60_combout ),
	.cout());
defparam \ram_in_reg[7][9]~60 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][9]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][9]~62 (
	.dataa(tdl_arr_9_11),
	.datab(reg_no_twiddle619),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][9]~62_combout ),
	.cout());
defparam \ram_in_reg[5][9]~62 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][9]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][9]~61 (
	.dataa(reg_no_twiddle619),
	.datab(tdl_arr_9_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][9]~61_combout ),
	.cout());
defparam \ram_in_reg[4][9]~61 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][9]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][9]~63 (
	.dataa(tdl_arr_9_13),
	.datab(tdl_arr_9_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][9]~63_combout ),
	.cout());
defparam \ram_in_reg[6][9]~63 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][9]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][8]~48 (
	.dataa(tdl_arr_8_14),
	.datab(tdl_arr_8_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][8]~48_combout ),
	.cout());
defparam \ram_in_reg[3][8]~48 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][8]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][8]~50 (
	.dataa(tdl_arr_8_1),
	.datab(reg_no_twiddle608),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][8]~50_combout ),
	.cout());
defparam \ram_in_reg[1][8]~50 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][8]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][8]~49 (
	.dataa(reg_no_twiddle608),
	.datab(tdl_arr_8_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][8]~49_combout ),
	.cout());
defparam \ram_in_reg[0][8]~49 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][8]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][8]~51 (
	.dataa(tdl_arr_8_12),
	.datab(tdl_arr_8_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][8]~51_combout ),
	.cout());
defparam \ram_in_reg[2][8]~51 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][8]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][8]~52 (
	.dataa(tdl_arr_8_15),
	.datab(tdl_arr_8_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][8]~52_combout ),
	.cout());
defparam \ram_in_reg[7][8]~52 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][8]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][8]~54 (
	.dataa(tdl_arr_8_11),
	.datab(reg_no_twiddle618),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][8]~54_combout ),
	.cout());
defparam \ram_in_reg[5][8]~54 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][8]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][8]~53 (
	.dataa(reg_no_twiddle618),
	.datab(tdl_arr_8_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][8]~53_combout ),
	.cout());
defparam \ram_in_reg[4][8]~53 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][8]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][8]~55 (
	.dataa(tdl_arr_8_13),
	.datab(tdl_arr_8_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][8]~55_combout ),
	.cout());
defparam \ram_in_reg[6][8]~55 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][8]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][7]~40 (
	.dataa(tdl_arr_7_14),
	.datab(tdl_arr_7_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~40_combout ),
	.cout());
defparam \ram_in_reg[3][7]~40 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][7]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][7]~42 (
	.dataa(tdl_arr_7_1),
	.datab(reg_no_twiddle607),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][7]~42_combout ),
	.cout());
defparam \ram_in_reg[1][7]~42 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][7]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][7]~41 (
	.dataa(reg_no_twiddle607),
	.datab(tdl_arr_7_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][7]~41_combout ),
	.cout());
defparam \ram_in_reg[0][7]~41 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][7]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][7]~43 (
	.dataa(tdl_arr_7_12),
	.datab(tdl_arr_7_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][7]~43_combout ),
	.cout());
defparam \ram_in_reg[2][7]~43 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][7]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][7]~44 (
	.dataa(tdl_arr_7_15),
	.datab(tdl_arr_7_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][7]~44_combout ),
	.cout());
defparam \ram_in_reg[7][7]~44 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][7]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][7]~46 (
	.dataa(tdl_arr_7_11),
	.datab(reg_no_twiddle617),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][7]~46_combout ),
	.cout());
defparam \ram_in_reg[5][7]~46 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][7]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][7]~45 (
	.dataa(reg_no_twiddle617),
	.datab(tdl_arr_7_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][7]~45_combout ),
	.cout());
defparam \ram_in_reg[4][7]~45 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][7]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][7]~47 (
	.dataa(tdl_arr_7_13),
	.datab(tdl_arr_7_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][7]~47_combout ),
	.cout());
defparam \ram_in_reg[6][7]~47 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][7]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][6]~32 (
	.dataa(tdl_arr_6_14),
	.datab(tdl_arr_6_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][6]~32_combout ),
	.cout());
defparam \ram_in_reg[3][6]~32 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][6]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][6]~34 (
	.dataa(tdl_arr_6_1),
	.datab(reg_no_twiddle606),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~34_combout ),
	.cout());
defparam \ram_in_reg[1][6]~34 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][6]~33 (
	.dataa(reg_no_twiddle606),
	.datab(tdl_arr_6_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][6]~33_combout ),
	.cout());
defparam \ram_in_reg[0][6]~33 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][6]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][6]~35 (
	.dataa(tdl_arr_6_12),
	.datab(tdl_arr_6_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][6]~35_combout ),
	.cout());
defparam \ram_in_reg[2][6]~35 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][6]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][6]~36 (
	.dataa(tdl_arr_6_15),
	.datab(tdl_arr_6_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][6]~36_combout ),
	.cout());
defparam \ram_in_reg[7][6]~36 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][6]~38 (
	.dataa(tdl_arr_6_11),
	.datab(reg_no_twiddle616),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][6]~38_combout ),
	.cout());
defparam \ram_in_reg[5][6]~38 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][6]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][6]~37 (
	.dataa(reg_no_twiddle616),
	.datab(tdl_arr_6_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][6]~37_combout ),
	.cout());
defparam \ram_in_reg[4][6]~37 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][6]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][6]~39 (
	.dataa(tdl_arr_6_13),
	.datab(tdl_arr_6_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][6]~39_combout ),
	.cout());
defparam \ram_in_reg[6][6]~39 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][6]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][5]~24 (
	.dataa(tdl_arr_5_14),
	.datab(tdl_arr_5_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~24_combout ),
	.cout());
defparam \ram_in_reg[3][5]~24 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][5]~26 (
	.dataa(tdl_arr_5_1),
	.datab(reg_no_twiddle605),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~26_combout ),
	.cout());
defparam \ram_in_reg[1][5]~26 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][5]~25 (
	.dataa(reg_no_twiddle605),
	.datab(tdl_arr_5_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~25_combout ),
	.cout());
defparam \ram_in_reg[0][5]~25 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][5]~27 (
	.dataa(tdl_arr_5_12),
	.datab(tdl_arr_5_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~27_combout ),
	.cout());
defparam \ram_in_reg[2][5]~27 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][5]~28 (
	.dataa(tdl_arr_5_15),
	.datab(tdl_arr_5_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][5]~28_combout ),
	.cout());
defparam \ram_in_reg[7][5]~28 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][5]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][5]~30 (
	.dataa(tdl_arr_5_11),
	.datab(reg_no_twiddle615),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][5]~30_combout ),
	.cout());
defparam \ram_in_reg[5][5]~30 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][5]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][5]~29 (
	.dataa(reg_no_twiddle615),
	.datab(tdl_arr_5_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][5]~29_combout ),
	.cout());
defparam \ram_in_reg[4][5]~29 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][5]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][5]~31 (
	.dataa(tdl_arr_5_13),
	.datab(tdl_arr_5_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][5]~31_combout ),
	.cout());
defparam \ram_in_reg[6][5]~31 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][5]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][4]~16 (
	.dataa(tdl_arr_4_1),
	.datab(tdl_arr_4_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][4]~16_combout ),
	.cout());
defparam \ram_in_reg[3][4]~16 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][4]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][4]~18 (
	.dataa(tdl_arr_4_12),
	.datab(reg_no_twiddle604),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][4]~18_combout ),
	.cout());
defparam \ram_in_reg[1][4]~18 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][4]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][4]~17 (
	.dataa(reg_no_twiddle604),
	.datab(tdl_arr_4_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][4]~17_combout ),
	.cout());
defparam \ram_in_reg[0][4]~17 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][4]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][4]~19 (
	.dataa(tdl_arr_4_11),
	.datab(tdl_arr_4_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][4]~19_combout ),
	.cout());
defparam \ram_in_reg[2][4]~19 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][4]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][4]~20 (
	.dataa(tdl_arr_4_13),
	.datab(tdl_arr_4_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][4]~20_combout ),
	.cout());
defparam \ram_in_reg[7][4]~20 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][4]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][4]~22 (
	.dataa(tdl_arr_4_15),
	.datab(reg_no_twiddle614),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][4]~22_combout ),
	.cout());
defparam \ram_in_reg[5][4]~22 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][4]~21 (
	.dataa(reg_no_twiddle614),
	.datab(tdl_arr_4_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][4]~21_combout ),
	.cout());
defparam \ram_in_reg[4][4]~21 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][4]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][4]~23 (
	.dataa(tdl_arr_4_14),
	.datab(tdl_arr_4_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][4]~23_combout ),
	.cout());
defparam \ram_in_reg[6][4]~23 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][4]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][3]~8 (
	.dataa(tdl_arr_3_1),
	.datab(tdl_arr_3_11),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~8_combout ),
	.cout());
defparam \ram_in_reg[3][3]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][3]~10 (
	.dataa(tdl_arr_3_12),
	.datab(reg_no_twiddle603),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~10_combout ),
	.cout());
defparam \ram_in_reg[1][3]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][3]~9 (
	.dataa(reg_no_twiddle603),
	.datab(tdl_arr_3_1),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~9_combout ),
	.cout());
defparam \ram_in_reg[0][3]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][3]~11 (
	.dataa(tdl_arr_3_11),
	.datab(tdl_arr_3_12),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~11_combout ),
	.cout());
defparam \ram_in_reg[2][3]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][3]~12 (
	.dataa(tdl_arr_3_13),
	.datab(tdl_arr_3_14),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[7][3]~12_combout ),
	.cout());
defparam \ram_in_reg[7][3]~12 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][3]~14 (
	.dataa(tdl_arr_3_15),
	.datab(reg_no_twiddle613),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[5][3]~14_combout ),
	.cout());
defparam \ram_in_reg[5][3]~14 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][3]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][3]~13 (
	.dataa(reg_no_twiddle613),
	.datab(tdl_arr_3_13),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[4][3]~13_combout ),
	.cout());
defparam \ram_in_reg[4][3]~13 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][3]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][3]~15 (
	.dataa(tdl_arr_3_14),
	.datab(tdl_arr_3_15),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_in_reg[6][3]~15_combout ),
	.cout());
defparam \ram_in_reg[6][3]~15 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][3]~15 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_data_r (
	ram_in_reg_2_3,
	ram_in_reg_2_7,
	ram_in_reg_2_1,
	ram_in_reg_2_5,
	ram_in_reg_1_3,
	ram_in_reg_1_7,
	ram_in_reg_1_1,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	ram_in_reg_0_1,
	ram_in_reg_0_5,
	ram_in_reg_2_6,
	ram_in_reg_2_4,
	ram_in_reg_1_6,
	ram_in_reg_1_4,
	ram_in_reg_0_6,
	ram_in_reg_0_4,
	ram_in_reg_9_3,
	ram_in_reg_9_7,
	ram_in_reg_9_1,
	ram_in_reg_9_5,
	ram_in_reg_8_3,
	ram_in_reg_8_7,
	ram_in_reg_8_1,
	ram_in_reg_8_5,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_9_6,
	ram_in_reg_9_4,
	ram_in_reg_8_6,
	ram_in_reg_8_4,
	ram_in_reg_7_6,
	ram_in_reg_7_4,
	ram_in_reg_6_6,
	ram_in_reg_6_4,
	ram_in_reg_5_6,
	ram_in_reg_5_4,
	ram_in_reg_4_6,
	ram_in_reg_4_4,
	ram_in_reg_3_6,
	ram_in_reg_3_4,
	ram_in_reg_2_2,
	ram_in_reg_2_0,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	ram_in_reg_0_2,
	ram_in_reg_0_0,
	ram_in_reg_9_2,
	ram_in_reg_9_0,
	ram_in_reg_8_2,
	ram_in_reg_8_0,
	ram_in_reg_7_2,
	ram_in_reg_7_0,
	ram_in_reg_6_2,
	ram_in_reg_6_0,
	ram_in_reg_5_2,
	ram_in_reg_5_0,
	ram_in_reg_4_2,
	ram_in_reg_4_0,
	ram_in_reg_3_2,
	ram_in_reg_3_0,
	global_clock_enable,
	lpp_ram_data_out_12_3,
	lpp_ram_data_out_12_0,
	tdl_arr_0_4,
	lpp_ram_data_out_12_1,
	lpp_ram_data_out_12_2,
	tdl_arr_1_4,
	lpp_ram_data_out_2_3,
	lpp_ram_data_out_2_0,
	lpp_ram_data_out_2_1,
	lpp_ram_data_out_2_2,
	lpp_ram_data_out_11_3,
	lpp_ram_data_out_11_0,
	lpp_ram_data_out_11_1,
	lpp_ram_data_out_11_2,
	lpp_ram_data_out_1_3,
	lpp_ram_data_out_1_0,
	lpp_ram_data_out_1_1,
	lpp_ram_data_out_1_2,
	lpp_ram_data_out_10_3,
	lpp_ram_data_out_10_0,
	lpp_ram_data_out_10_1,
	lpp_ram_data_out_10_2,
	lpp_ram_data_out_0_3,
	lpp_ram_data_out_0_0,
	lpp_ram_data_out_0_1,
	lpp_ram_data_out_0_2,
	lpp_ram_data_out_19_3,
	lpp_ram_data_out_19_0,
	lpp_ram_data_out_19_1,
	lpp_ram_data_out_19_2,
	lpp_ram_data_out_9_3,
	lpp_ram_data_out_9_0,
	lpp_ram_data_out_9_1,
	lpp_ram_data_out_9_2,
	lpp_ram_data_out_18_3,
	lpp_ram_data_out_18_0,
	lpp_ram_data_out_18_1,
	lpp_ram_data_out_18_2,
	lpp_ram_data_out_8_3,
	lpp_ram_data_out_8_0,
	lpp_ram_data_out_8_1,
	lpp_ram_data_out_8_2,
	lpp_ram_data_out_17_3,
	lpp_ram_data_out_17_0,
	lpp_ram_data_out_17_1,
	lpp_ram_data_out_17_2,
	lpp_ram_data_out_7_3,
	lpp_ram_data_out_7_0,
	lpp_ram_data_out_7_1,
	lpp_ram_data_out_7_2,
	lpp_ram_data_out_16_3,
	lpp_ram_data_out_16_0,
	lpp_ram_data_out_16_1,
	lpp_ram_data_out_16_2,
	lpp_ram_data_out_6_3,
	lpp_ram_data_out_6_0,
	lpp_ram_data_out_6_1,
	lpp_ram_data_out_6_2,
	lpp_ram_data_out_15_3,
	lpp_ram_data_out_15_0,
	lpp_ram_data_out_15_1,
	lpp_ram_data_out_15_2,
	lpp_ram_data_out_5_3,
	lpp_ram_data_out_5_0,
	lpp_ram_data_out_5_1,
	lpp_ram_data_out_5_2,
	lpp_ram_data_out_14_3,
	lpp_ram_data_out_14_0,
	lpp_ram_data_out_14_1,
	lpp_ram_data_out_14_2,
	lpp_ram_data_out_4_3,
	lpp_ram_data_out_4_0,
	lpp_ram_data_out_4_1,
	lpp_ram_data_out_4_2,
	lpp_ram_data_out_13_3,
	lpp_ram_data_out_13_0,
	lpp_ram_data_out_13_1,
	lpp_ram_data_out_13_2,
	lpp_ram_data_out_3_3,
	lpp_ram_data_out_3_0,
	lpp_ram_data_out_3_1,
	lpp_ram_data_out_3_2,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_2_3;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_1;
output 	ram_in_reg_2_5;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_7;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_5;
output 	ram_in_reg_0_3;
output 	ram_in_reg_0_7;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_5;
output 	ram_in_reg_2_6;
output 	ram_in_reg_2_4;
output 	ram_in_reg_1_6;
output 	ram_in_reg_1_4;
output 	ram_in_reg_0_6;
output 	ram_in_reg_0_4;
output 	ram_in_reg_9_3;
output 	ram_in_reg_9_7;
output 	ram_in_reg_9_1;
output 	ram_in_reg_9_5;
output 	ram_in_reg_8_3;
output 	ram_in_reg_8_7;
output 	ram_in_reg_8_1;
output 	ram_in_reg_8_5;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_7;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_5;
output 	ram_in_reg_6_3;
output 	ram_in_reg_6_7;
output 	ram_in_reg_6_1;
output 	ram_in_reg_6_5;
output 	ram_in_reg_5_3;
output 	ram_in_reg_5_7;
output 	ram_in_reg_5_1;
output 	ram_in_reg_5_5;
output 	ram_in_reg_4_3;
output 	ram_in_reg_4_7;
output 	ram_in_reg_4_1;
output 	ram_in_reg_4_5;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_7;
output 	ram_in_reg_3_1;
output 	ram_in_reg_3_5;
output 	ram_in_reg_9_6;
output 	ram_in_reg_9_4;
output 	ram_in_reg_8_6;
output 	ram_in_reg_8_4;
output 	ram_in_reg_7_6;
output 	ram_in_reg_7_4;
output 	ram_in_reg_6_6;
output 	ram_in_reg_6_4;
output 	ram_in_reg_5_6;
output 	ram_in_reg_5_4;
output 	ram_in_reg_4_6;
output 	ram_in_reg_4_4;
output 	ram_in_reg_3_6;
output 	ram_in_reg_3_4;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_0;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_0;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_0;
output 	ram_in_reg_9_2;
output 	ram_in_reg_9_0;
output 	ram_in_reg_8_2;
output 	ram_in_reg_8_0;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_0;
output 	ram_in_reg_6_2;
output 	ram_in_reg_6_0;
output 	ram_in_reg_5_2;
output 	ram_in_reg_5_0;
output 	ram_in_reg_4_2;
output 	ram_in_reg_4_0;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_0;
input 	global_clock_enable;
input 	lpp_ram_data_out_12_3;
input 	lpp_ram_data_out_12_0;
input 	tdl_arr_0_4;
input 	lpp_ram_data_out_12_1;
input 	lpp_ram_data_out_12_2;
input 	tdl_arr_1_4;
input 	lpp_ram_data_out_2_3;
input 	lpp_ram_data_out_2_0;
input 	lpp_ram_data_out_2_1;
input 	lpp_ram_data_out_2_2;
input 	lpp_ram_data_out_11_3;
input 	lpp_ram_data_out_11_0;
input 	lpp_ram_data_out_11_1;
input 	lpp_ram_data_out_11_2;
input 	lpp_ram_data_out_1_3;
input 	lpp_ram_data_out_1_0;
input 	lpp_ram_data_out_1_1;
input 	lpp_ram_data_out_1_2;
input 	lpp_ram_data_out_10_3;
input 	lpp_ram_data_out_10_0;
input 	lpp_ram_data_out_10_1;
input 	lpp_ram_data_out_10_2;
input 	lpp_ram_data_out_0_3;
input 	lpp_ram_data_out_0_0;
input 	lpp_ram_data_out_0_1;
input 	lpp_ram_data_out_0_2;
input 	lpp_ram_data_out_19_3;
input 	lpp_ram_data_out_19_0;
input 	lpp_ram_data_out_19_1;
input 	lpp_ram_data_out_19_2;
input 	lpp_ram_data_out_9_3;
input 	lpp_ram_data_out_9_0;
input 	lpp_ram_data_out_9_1;
input 	lpp_ram_data_out_9_2;
input 	lpp_ram_data_out_18_3;
input 	lpp_ram_data_out_18_0;
input 	lpp_ram_data_out_18_1;
input 	lpp_ram_data_out_18_2;
input 	lpp_ram_data_out_8_3;
input 	lpp_ram_data_out_8_0;
input 	lpp_ram_data_out_8_1;
input 	lpp_ram_data_out_8_2;
input 	lpp_ram_data_out_17_3;
input 	lpp_ram_data_out_17_0;
input 	lpp_ram_data_out_17_1;
input 	lpp_ram_data_out_17_2;
input 	lpp_ram_data_out_7_3;
input 	lpp_ram_data_out_7_0;
input 	lpp_ram_data_out_7_1;
input 	lpp_ram_data_out_7_2;
input 	lpp_ram_data_out_16_3;
input 	lpp_ram_data_out_16_0;
input 	lpp_ram_data_out_16_1;
input 	lpp_ram_data_out_16_2;
input 	lpp_ram_data_out_6_3;
input 	lpp_ram_data_out_6_0;
input 	lpp_ram_data_out_6_1;
input 	lpp_ram_data_out_6_2;
input 	lpp_ram_data_out_15_3;
input 	lpp_ram_data_out_15_0;
input 	lpp_ram_data_out_15_1;
input 	lpp_ram_data_out_15_2;
input 	lpp_ram_data_out_5_3;
input 	lpp_ram_data_out_5_0;
input 	lpp_ram_data_out_5_1;
input 	lpp_ram_data_out_5_2;
input 	lpp_ram_data_out_14_3;
input 	lpp_ram_data_out_14_0;
input 	lpp_ram_data_out_14_1;
input 	lpp_ram_data_out_14_2;
input 	lpp_ram_data_out_4_3;
input 	lpp_ram_data_out_4_0;
input 	lpp_ram_data_out_4_1;
input 	lpp_ram_data_out_4_2;
input 	lpp_ram_data_out_13_3;
input 	lpp_ram_data_out_13_0;
input 	lpp_ram_data_out_13_1;
input 	lpp_ram_data_out_13_2;
input 	lpp_ram_data_out_3_3;
input 	lpp_ram_data_out_3_0;
input 	lpp_ram_data_out_3_1;
input 	lpp_ram_data_out_3_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[3][2]~0_combout ;
wire \ram_in_reg[1][2]~2_combout ;
wire \ram_in_reg[7][2]~1_combout ;
wire \ram_in_reg[5][2]~3_combout ;
wire \ram_in_reg[3][1]~64_combout ;
wire \ram_in_reg[1][1]~66_combout ;
wire \ram_in_reg[7][1]~65_combout ;
wire \ram_in_reg[5][1]~67_combout ;
wire \ram_in_reg[3][0]~72_combout ;
wire \ram_in_reg[1][0]~74_combout ;
wire \ram_in_reg[7][0]~73_combout ;
wire \ram_in_reg[5][0]~75_combout ;
wire \ram_in_reg[6][2]~6_combout ;
wire \ram_in_reg[4][2]~7_combout ;
wire \ram_in_reg[6][1]~70_combout ;
wire \ram_in_reg[4][1]~71_combout ;
wire \ram_in_reg[6][0]~78_combout ;
wire \ram_in_reg[4][0]~79_combout ;
wire \ram_in_reg[3][9]~56_combout ;
wire \ram_in_reg[1][9]~58_combout ;
wire \ram_in_reg[7][9]~57_combout ;
wire \ram_in_reg[5][9]~59_combout ;
wire \ram_in_reg[3][8]~48_combout ;
wire \ram_in_reg[1][8]~50_combout ;
wire \ram_in_reg[7][8]~49_combout ;
wire \ram_in_reg[5][8]~51_combout ;
wire \ram_in_reg[3][7]~40_combout ;
wire \ram_in_reg[1][7]~42_combout ;
wire \ram_in_reg[7][7]~41_combout ;
wire \ram_in_reg[5][7]~43_combout ;
wire \ram_in_reg[3][6]~32_combout ;
wire \ram_in_reg[1][6]~34_combout ;
wire \ram_in_reg[7][6]~33_combout ;
wire \ram_in_reg[5][6]~35_combout ;
wire \ram_in_reg[3][5]~24_combout ;
wire \ram_in_reg[1][5]~26_combout ;
wire \ram_in_reg[7][5]~25_combout ;
wire \ram_in_reg[5][5]~27_combout ;
wire \ram_in_reg[3][4]~16_combout ;
wire \ram_in_reg[1][4]~18_combout ;
wire \ram_in_reg[7][4]~17_combout ;
wire \ram_in_reg[5][4]~19_combout ;
wire \ram_in_reg[3][3]~8_combout ;
wire \ram_in_reg[1][3]~10_combout ;
wire \ram_in_reg[7][3]~9_combout ;
wire \ram_in_reg[5][3]~11_combout ;
wire \ram_in_reg[6][9]~62_combout ;
wire \ram_in_reg[4][9]~63_combout ;
wire \ram_in_reg[6][8]~54_combout ;
wire \ram_in_reg[4][8]~55_combout ;
wire \ram_in_reg[6][7]~46_combout ;
wire \ram_in_reg[4][7]~47_combout ;
wire \ram_in_reg[6][6]~38_combout ;
wire \ram_in_reg[4][6]~39_combout ;
wire \ram_in_reg[6][5]~30_combout ;
wire \ram_in_reg[4][5]~31_combout ;
wire \ram_in_reg[6][4]~22_combout ;
wire \ram_in_reg[4][4]~23_combout ;
wire \ram_in_reg[6][3]~14_combout ;
wire \ram_in_reg[4][3]~15_combout ;
wire \ram_in_reg[2][2]~4_combout ;
wire \ram_in_reg[0][2]~5_combout ;
wire \ram_in_reg[2][1]~68_combout ;
wire \ram_in_reg[0][1]~69_combout ;
wire \ram_in_reg[2][0]~76_combout ;
wire \ram_in_reg[0][0]~77_combout ;
wire \ram_in_reg[2][9]~60_combout ;
wire \ram_in_reg[0][9]~61_combout ;
wire \ram_in_reg[2][8]~52_combout ;
wire \ram_in_reg[0][8]~53_combout ;
wire \ram_in_reg[2][7]~44_combout ;
wire \ram_in_reg[0][7]~45_combout ;
wire \ram_in_reg[2][6]~36_combout ;
wire \ram_in_reg[0][6]~37_combout ;
wire \ram_in_reg[2][5]~28_combout ;
wire \ram_in_reg[0][5]~29_combout ;
wire \ram_in_reg[2][4]~20_combout ;
wire \ram_in_reg[0][4]~21_combout ;
wire \ram_in_reg[2][3]~12_combout ;
wire \ram_in_reg[0][3]~13_combout ;


dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\ram_in_reg[3][2]~0_combout ),
	.asdata(\ram_in_reg[1][2]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\ram_in_reg[7][2]~1_combout ),
	.asdata(\ram_in_reg[5][2]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~2_combout ),
	.asdata(\ram_in_reg[3][2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\ram_in_reg[5][2]~3_combout ),
	.asdata(\ram_in_reg[7][2]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~64_combout ),
	.asdata(\ram_in_reg[1][1]~66_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\ram_in_reg[7][1]~65_combout ),
	.asdata(\ram_in_reg[5][1]~67_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~66_combout ),
	.asdata(\ram_in_reg[3][1]~64_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\ram_in_reg[5][1]~67_combout ),
	.asdata(\ram_in_reg[7][1]~65_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\ram_in_reg[3][0]~72_combout ),
	.asdata(\ram_in_reg[1][0]~74_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\ram_in_reg[7][0]~73_combout ),
	.asdata(\ram_in_reg[5][0]~75_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\ram_in_reg[1][0]~74_combout ),
	.asdata(\ram_in_reg[3][0]~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\ram_in_reg[5][0]~75_combout ),
	.asdata(\ram_in_reg[7][0]~73_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\ram_in_reg[6][2]~6_combout ),
	.asdata(\ram_in_reg[4][2]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\ram_in_reg[4][2]~7_combout ),
	.asdata(\ram_in_reg[6][2]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\ram_in_reg[6][1]~70_combout ),
	.asdata(\ram_in_reg[4][1]~71_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\ram_in_reg[4][1]~71_combout ),
	.asdata(\ram_in_reg[6][1]~70_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\ram_in_reg[6][0]~78_combout ),
	.asdata(\ram_in_reg[4][0]~79_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\ram_in_reg[4][0]~79_combout ),
	.asdata(\ram_in_reg[6][0]~78_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[3][9] (
	.clk(clk),
	.d(\ram_in_reg[3][9]~56_combout ),
	.asdata(\ram_in_reg[1][9]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_3),
	.prn(vcc));
defparam \ram_in_reg[3][9] .is_wysiwyg = "true";
defparam \ram_in_reg[3][9] .power_up = "low";

dffeas \ram_in_reg[7][9] (
	.clk(clk),
	.d(\ram_in_reg[7][9]~57_combout ),
	.asdata(\ram_in_reg[5][9]~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_7),
	.prn(vcc));
defparam \ram_in_reg[7][9] .is_wysiwyg = "true";
defparam \ram_in_reg[7][9] .power_up = "low";

dffeas \ram_in_reg[1][9] (
	.clk(clk),
	.d(\ram_in_reg[1][9]~58_combout ),
	.asdata(\ram_in_reg[3][9]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_1),
	.prn(vcc));
defparam \ram_in_reg[1][9] .is_wysiwyg = "true";
defparam \ram_in_reg[1][9] .power_up = "low";

dffeas \ram_in_reg[5][9] (
	.clk(clk),
	.d(\ram_in_reg[5][9]~59_combout ),
	.asdata(\ram_in_reg[7][9]~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_5),
	.prn(vcc));
defparam \ram_in_reg[5][9] .is_wysiwyg = "true";
defparam \ram_in_reg[5][9] .power_up = "low";

dffeas \ram_in_reg[3][8] (
	.clk(clk),
	.d(\ram_in_reg[3][8]~48_combout ),
	.asdata(\ram_in_reg[1][8]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_3),
	.prn(vcc));
defparam \ram_in_reg[3][8] .is_wysiwyg = "true";
defparam \ram_in_reg[3][8] .power_up = "low";

dffeas \ram_in_reg[7][8] (
	.clk(clk),
	.d(\ram_in_reg[7][8]~49_combout ),
	.asdata(\ram_in_reg[5][8]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_7),
	.prn(vcc));
defparam \ram_in_reg[7][8] .is_wysiwyg = "true";
defparam \ram_in_reg[7][8] .power_up = "low";

dffeas \ram_in_reg[1][8] (
	.clk(clk),
	.d(\ram_in_reg[1][8]~50_combout ),
	.asdata(\ram_in_reg[3][8]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_1),
	.prn(vcc));
defparam \ram_in_reg[1][8] .is_wysiwyg = "true";
defparam \ram_in_reg[1][8] .power_up = "low";

dffeas \ram_in_reg[5][8] (
	.clk(clk),
	.d(\ram_in_reg[5][8]~51_combout ),
	.asdata(\ram_in_reg[7][8]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_5),
	.prn(vcc));
defparam \ram_in_reg[5][8] .is_wysiwyg = "true";
defparam \ram_in_reg[5][8] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~40_combout ),
	.asdata(\ram_in_reg[1][7]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\ram_in_reg[7][7]~41_combout ),
	.asdata(\ram_in_reg[5][7]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\ram_in_reg[1][7]~42_combout ),
	.asdata(\ram_in_reg[3][7]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\ram_in_reg[5][7]~43_combout ),
	.asdata(\ram_in_reg[7][7]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\ram_in_reg[3][6]~32_combout ),
	.asdata(\ram_in_reg[1][6]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\ram_in_reg[7][6]~33_combout ),
	.asdata(\ram_in_reg[5][6]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~34_combout ),
	.asdata(\ram_in_reg[3][6]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\ram_in_reg[5][6]~35_combout ),
	.asdata(\ram_in_reg[7][6]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~24_combout ),
	.asdata(\ram_in_reg[1][5]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\ram_in_reg[7][5]~25_combout ),
	.asdata(\ram_in_reg[5][5]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~26_combout ),
	.asdata(\ram_in_reg[3][5]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\ram_in_reg[5][5]~27_combout ),
	.asdata(\ram_in_reg[7][5]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\ram_in_reg[3][4]~16_combout ),
	.asdata(\ram_in_reg[1][4]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\ram_in_reg[7][4]~17_combout ),
	.asdata(\ram_in_reg[5][4]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\ram_in_reg[1][4]~18_combout ),
	.asdata(\ram_in_reg[3][4]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\ram_in_reg[5][4]~19_combout ),
	.asdata(\ram_in_reg[7][4]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~8_combout ),
	.asdata(\ram_in_reg[1][3]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\ram_in_reg[7][3]~9_combout ),
	.asdata(\ram_in_reg[5][3]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~10_combout ),
	.asdata(\ram_in_reg[3][3]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\ram_in_reg[5][3]~11_combout ),
	.asdata(\ram_in_reg[7][3]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[6][9] (
	.clk(clk),
	.d(\ram_in_reg[6][9]~62_combout ),
	.asdata(\ram_in_reg[4][9]~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_6),
	.prn(vcc));
defparam \ram_in_reg[6][9] .is_wysiwyg = "true";
defparam \ram_in_reg[6][9] .power_up = "low";

dffeas \ram_in_reg[4][9] (
	.clk(clk),
	.d(\ram_in_reg[4][9]~63_combout ),
	.asdata(\ram_in_reg[6][9]~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_4),
	.prn(vcc));
defparam \ram_in_reg[4][9] .is_wysiwyg = "true";
defparam \ram_in_reg[4][9] .power_up = "low";

dffeas \ram_in_reg[6][8] (
	.clk(clk),
	.d(\ram_in_reg[6][8]~54_combout ),
	.asdata(\ram_in_reg[4][8]~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_6),
	.prn(vcc));
defparam \ram_in_reg[6][8] .is_wysiwyg = "true";
defparam \ram_in_reg[6][8] .power_up = "low";

dffeas \ram_in_reg[4][8] (
	.clk(clk),
	.d(\ram_in_reg[4][8]~55_combout ),
	.asdata(\ram_in_reg[6][8]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_4),
	.prn(vcc));
defparam \ram_in_reg[4][8] .is_wysiwyg = "true";
defparam \ram_in_reg[4][8] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\ram_in_reg[6][7]~46_combout ),
	.asdata(\ram_in_reg[4][7]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\ram_in_reg[4][7]~47_combout ),
	.asdata(\ram_in_reg[6][7]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\ram_in_reg[6][6]~38_combout ),
	.asdata(\ram_in_reg[4][6]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\ram_in_reg[4][6]~39_combout ),
	.asdata(\ram_in_reg[6][6]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\ram_in_reg[6][5]~30_combout ),
	.asdata(\ram_in_reg[4][5]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\ram_in_reg[4][5]~31_combout ),
	.asdata(\ram_in_reg[6][5]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\ram_in_reg[6][4]~22_combout ),
	.asdata(\ram_in_reg[4][4]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\ram_in_reg[4][4]~23_combout ),
	.asdata(\ram_in_reg[6][4]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\ram_in_reg[6][3]~14_combout ),
	.asdata(\ram_in_reg[4][3]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\ram_in_reg[4][3]~15_combout ),
	.asdata(\ram_in_reg[6][3]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\ram_in_reg[2][2]~4_combout ),
	.asdata(\ram_in_reg[0][2]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\ram_in_reg[0][2]~5_combout ),
	.asdata(\ram_in_reg[2][2]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~68_combout ),
	.asdata(\ram_in_reg[0][1]~69_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~69_combout ),
	.asdata(\ram_in_reg[2][1]~68_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\ram_in_reg[2][0]~76_combout ),
	.asdata(\ram_in_reg[0][0]~77_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\ram_in_reg[0][0]~77_combout ),
	.asdata(\ram_in_reg[2][0]~76_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[2][9] (
	.clk(clk),
	.d(\ram_in_reg[2][9]~60_combout ),
	.asdata(\ram_in_reg[0][9]~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_2),
	.prn(vcc));
defparam \ram_in_reg[2][9] .is_wysiwyg = "true";
defparam \ram_in_reg[2][9] .power_up = "low";

dffeas \ram_in_reg[0][9] (
	.clk(clk),
	.d(\ram_in_reg[0][9]~61_combout ),
	.asdata(\ram_in_reg[2][9]~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_0),
	.prn(vcc));
defparam \ram_in_reg[0][9] .is_wysiwyg = "true";
defparam \ram_in_reg[0][9] .power_up = "low";

dffeas \ram_in_reg[2][8] (
	.clk(clk),
	.d(\ram_in_reg[2][8]~52_combout ),
	.asdata(\ram_in_reg[0][8]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_2),
	.prn(vcc));
defparam \ram_in_reg[2][8] .is_wysiwyg = "true";
defparam \ram_in_reg[2][8] .power_up = "low";

dffeas \ram_in_reg[0][8] (
	.clk(clk),
	.d(\ram_in_reg[0][8]~53_combout ),
	.asdata(\ram_in_reg[2][8]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_0),
	.prn(vcc));
defparam \ram_in_reg[0][8] .is_wysiwyg = "true";
defparam \ram_in_reg[0][8] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\ram_in_reg[2][7]~44_combout ),
	.asdata(\ram_in_reg[0][7]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\ram_in_reg[0][7]~45_combout ),
	.asdata(\ram_in_reg[2][7]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\ram_in_reg[2][6]~36_combout ),
	.asdata(\ram_in_reg[0][6]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\ram_in_reg[0][6]~37_combout ),
	.asdata(\ram_in_reg[2][6]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~28_combout ),
	.asdata(\ram_in_reg[0][5]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~29_combout ),
	.asdata(\ram_in_reg[2][5]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\ram_in_reg[2][4]~20_combout ),
	.asdata(\ram_in_reg[0][4]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\ram_in_reg[0][4]~21_combout ),
	.asdata(\ram_in_reg[2][4]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~12_combout ),
	.asdata(\ram_in_reg[0][3]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~13_combout ),
	.asdata(\ram_in_reg[2][3]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(tdl_arr_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

cycloneive_lcell_comb \ram_in_reg[3][2]~0 (
	.dataa(lpp_ram_data_out_12_3),
	.datab(lpp_ram_data_out_12_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][2]~0_combout ),
	.cout());
defparam \ram_in_reg[3][2]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][2]~2 (
	.dataa(lpp_ram_data_out_12_1),
	.datab(lpp_ram_data_out_12_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][2]~2_combout ),
	.cout());
defparam \ram_in_reg[1][2]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][2]~1 (
	.dataa(lpp_ram_data_out_2_3),
	.datab(lpp_ram_data_out_2_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][2]~1_combout ),
	.cout());
defparam \ram_in_reg[7][2]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][2]~3 (
	.dataa(lpp_ram_data_out_2_1),
	.datab(lpp_ram_data_out_2_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][2]~3_combout ),
	.cout());
defparam \ram_in_reg[5][2]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][1]~64 (
	.dataa(lpp_ram_data_out_11_3),
	.datab(lpp_ram_data_out_11_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~64_combout ),
	.cout());
defparam \ram_in_reg[3][1]~64 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][1]~66 (
	.dataa(lpp_ram_data_out_11_1),
	.datab(lpp_ram_data_out_11_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~66_combout ),
	.cout());
defparam \ram_in_reg[1][1]~66 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][1]~65 (
	.dataa(lpp_ram_data_out_1_3),
	.datab(lpp_ram_data_out_1_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][1]~65_combout ),
	.cout());
defparam \ram_in_reg[7][1]~65 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][1]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][1]~67 (
	.dataa(lpp_ram_data_out_1_1),
	.datab(lpp_ram_data_out_1_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][1]~67_combout ),
	.cout());
defparam \ram_in_reg[5][1]~67 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][1]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][0]~72 (
	.dataa(lpp_ram_data_out_10_3),
	.datab(lpp_ram_data_out_10_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][0]~72_combout ),
	.cout());
defparam \ram_in_reg[3][0]~72 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][0]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][0]~74 (
	.dataa(lpp_ram_data_out_10_1),
	.datab(lpp_ram_data_out_10_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][0]~74_combout ),
	.cout());
defparam \ram_in_reg[1][0]~74 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][0]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][0]~73 (
	.dataa(lpp_ram_data_out_0_3),
	.datab(lpp_ram_data_out_0_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][0]~73_combout ),
	.cout());
defparam \ram_in_reg[7][0]~73 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][0]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][0]~75 (
	.dataa(lpp_ram_data_out_0_1),
	.datab(lpp_ram_data_out_0_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][0]~75_combout ),
	.cout());
defparam \ram_in_reg[5][0]~75 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][0]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][2]~6 (
	.dataa(lpp_ram_data_out_2_2),
	.datab(lpp_ram_data_out_2_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][2]~6_combout ),
	.cout());
defparam \ram_in_reg[6][2]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][2]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][2]~7 (
	.dataa(lpp_ram_data_out_2_0),
	.datab(lpp_ram_data_out_2_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][2]~7_combout ),
	.cout());
defparam \ram_in_reg[4][2]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][2]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][1]~70 (
	.dataa(lpp_ram_data_out_1_2),
	.datab(lpp_ram_data_out_1_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][1]~70_combout ),
	.cout());
defparam \ram_in_reg[6][1]~70 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][1]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][1]~71 (
	.dataa(lpp_ram_data_out_1_0),
	.datab(lpp_ram_data_out_1_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][1]~71_combout ),
	.cout());
defparam \ram_in_reg[4][1]~71 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][1]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][0]~78 (
	.dataa(lpp_ram_data_out_0_2),
	.datab(lpp_ram_data_out_0_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][0]~78_combout ),
	.cout());
defparam \ram_in_reg[6][0]~78 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][0]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][0]~79 (
	.dataa(lpp_ram_data_out_0_0),
	.datab(lpp_ram_data_out_0_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][0]~79_combout ),
	.cout());
defparam \ram_in_reg[4][0]~79 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][0]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][9]~56 (
	.dataa(lpp_ram_data_out_19_3),
	.datab(lpp_ram_data_out_19_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][9]~56_combout ),
	.cout());
defparam \ram_in_reg[3][9]~56 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][9]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][9]~58 (
	.dataa(lpp_ram_data_out_19_1),
	.datab(lpp_ram_data_out_19_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][9]~58_combout ),
	.cout());
defparam \ram_in_reg[1][9]~58 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][9]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][9]~57 (
	.dataa(lpp_ram_data_out_9_3),
	.datab(lpp_ram_data_out_9_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][9]~57_combout ),
	.cout());
defparam \ram_in_reg[7][9]~57 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][9]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][9]~59 (
	.dataa(lpp_ram_data_out_9_1),
	.datab(lpp_ram_data_out_9_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][9]~59_combout ),
	.cout());
defparam \ram_in_reg[5][9]~59 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][9]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][8]~48 (
	.dataa(lpp_ram_data_out_18_3),
	.datab(lpp_ram_data_out_18_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][8]~48_combout ),
	.cout());
defparam \ram_in_reg[3][8]~48 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][8]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][8]~50 (
	.dataa(lpp_ram_data_out_18_1),
	.datab(lpp_ram_data_out_18_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][8]~50_combout ),
	.cout());
defparam \ram_in_reg[1][8]~50 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][8]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][8]~49 (
	.dataa(lpp_ram_data_out_8_3),
	.datab(lpp_ram_data_out_8_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][8]~49_combout ),
	.cout());
defparam \ram_in_reg[7][8]~49 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][8]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][8]~51 (
	.dataa(lpp_ram_data_out_8_1),
	.datab(lpp_ram_data_out_8_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][8]~51_combout ),
	.cout());
defparam \ram_in_reg[5][8]~51 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][8]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][7]~40 (
	.dataa(lpp_ram_data_out_17_3),
	.datab(lpp_ram_data_out_17_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~40_combout ),
	.cout());
defparam \ram_in_reg[3][7]~40 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][7]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][7]~42 (
	.dataa(lpp_ram_data_out_17_1),
	.datab(lpp_ram_data_out_17_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][7]~42_combout ),
	.cout());
defparam \ram_in_reg[1][7]~42 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][7]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][7]~41 (
	.dataa(lpp_ram_data_out_7_3),
	.datab(lpp_ram_data_out_7_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][7]~41_combout ),
	.cout());
defparam \ram_in_reg[7][7]~41 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][7]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][7]~43 (
	.dataa(lpp_ram_data_out_7_1),
	.datab(lpp_ram_data_out_7_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][7]~43_combout ),
	.cout());
defparam \ram_in_reg[5][7]~43 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][7]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][6]~32 (
	.dataa(lpp_ram_data_out_16_3),
	.datab(lpp_ram_data_out_16_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][6]~32_combout ),
	.cout());
defparam \ram_in_reg[3][6]~32 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][6]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][6]~34 (
	.dataa(lpp_ram_data_out_16_1),
	.datab(lpp_ram_data_out_16_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~34_combout ),
	.cout());
defparam \ram_in_reg[1][6]~34 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][6]~33 (
	.dataa(lpp_ram_data_out_6_3),
	.datab(lpp_ram_data_out_6_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][6]~33_combout ),
	.cout());
defparam \ram_in_reg[7][6]~33 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][6]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][6]~35 (
	.dataa(lpp_ram_data_out_6_1),
	.datab(lpp_ram_data_out_6_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][6]~35_combout ),
	.cout());
defparam \ram_in_reg[5][6]~35 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][6]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][5]~24 (
	.dataa(lpp_ram_data_out_15_3),
	.datab(lpp_ram_data_out_15_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~24_combout ),
	.cout());
defparam \ram_in_reg[3][5]~24 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][5]~26 (
	.dataa(lpp_ram_data_out_15_1),
	.datab(lpp_ram_data_out_15_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~26_combout ),
	.cout());
defparam \ram_in_reg[1][5]~26 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][5]~25 (
	.dataa(lpp_ram_data_out_5_3),
	.datab(lpp_ram_data_out_5_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][5]~25_combout ),
	.cout());
defparam \ram_in_reg[7][5]~25 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][5]~27 (
	.dataa(lpp_ram_data_out_5_1),
	.datab(lpp_ram_data_out_5_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][5]~27_combout ),
	.cout());
defparam \ram_in_reg[5][5]~27 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][5]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][4]~16 (
	.dataa(lpp_ram_data_out_14_3),
	.datab(lpp_ram_data_out_14_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][4]~16_combout ),
	.cout());
defparam \ram_in_reg[3][4]~16 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][4]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][4]~18 (
	.dataa(lpp_ram_data_out_14_1),
	.datab(lpp_ram_data_out_14_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][4]~18_combout ),
	.cout());
defparam \ram_in_reg[1][4]~18 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][4]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][4]~17 (
	.dataa(lpp_ram_data_out_4_3),
	.datab(lpp_ram_data_out_4_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][4]~17_combout ),
	.cout());
defparam \ram_in_reg[7][4]~17 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][4]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][4]~19 (
	.dataa(lpp_ram_data_out_4_1),
	.datab(lpp_ram_data_out_4_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][4]~19_combout ),
	.cout());
defparam \ram_in_reg[5][4]~19 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][4]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][3]~8 (
	.dataa(lpp_ram_data_out_13_3),
	.datab(lpp_ram_data_out_13_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~8_combout ),
	.cout());
defparam \ram_in_reg[3][3]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][3]~10 (
	.dataa(lpp_ram_data_out_13_1),
	.datab(lpp_ram_data_out_13_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~10_combout ),
	.cout());
defparam \ram_in_reg[1][3]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][3]~9 (
	.dataa(lpp_ram_data_out_3_3),
	.datab(lpp_ram_data_out_3_0),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][3]~9_combout ),
	.cout());
defparam \ram_in_reg[7][3]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][3]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][3]~11 (
	.dataa(lpp_ram_data_out_3_1),
	.datab(lpp_ram_data_out_3_2),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][3]~11_combout ),
	.cout());
defparam \ram_in_reg[5][3]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][3]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][9]~62 (
	.dataa(lpp_ram_data_out_9_2),
	.datab(lpp_ram_data_out_9_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][9]~62_combout ),
	.cout());
defparam \ram_in_reg[6][9]~62 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][9]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][9]~63 (
	.dataa(lpp_ram_data_out_9_0),
	.datab(lpp_ram_data_out_9_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][9]~63_combout ),
	.cout());
defparam \ram_in_reg[4][9]~63 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][9]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][8]~54 (
	.dataa(lpp_ram_data_out_8_2),
	.datab(lpp_ram_data_out_8_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][8]~54_combout ),
	.cout());
defparam \ram_in_reg[6][8]~54 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][8]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][8]~55 (
	.dataa(lpp_ram_data_out_8_0),
	.datab(lpp_ram_data_out_8_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][8]~55_combout ),
	.cout());
defparam \ram_in_reg[4][8]~55 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][8]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][7]~46 (
	.dataa(lpp_ram_data_out_7_2),
	.datab(lpp_ram_data_out_7_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][7]~46_combout ),
	.cout());
defparam \ram_in_reg[6][7]~46 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][7]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][7]~47 (
	.dataa(lpp_ram_data_out_7_0),
	.datab(lpp_ram_data_out_7_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][7]~47_combout ),
	.cout());
defparam \ram_in_reg[4][7]~47 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][7]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][6]~38 (
	.dataa(lpp_ram_data_out_6_2),
	.datab(lpp_ram_data_out_6_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][6]~38_combout ),
	.cout());
defparam \ram_in_reg[6][6]~38 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][6]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][6]~39 (
	.dataa(lpp_ram_data_out_6_0),
	.datab(lpp_ram_data_out_6_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][6]~39_combout ),
	.cout());
defparam \ram_in_reg[4][6]~39 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][6]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][5]~30 (
	.dataa(lpp_ram_data_out_5_2),
	.datab(lpp_ram_data_out_5_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][5]~30_combout ),
	.cout());
defparam \ram_in_reg[6][5]~30 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][5]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][5]~31 (
	.dataa(lpp_ram_data_out_5_0),
	.datab(lpp_ram_data_out_5_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][5]~31_combout ),
	.cout());
defparam \ram_in_reg[4][5]~31 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][5]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][4]~22 (
	.dataa(lpp_ram_data_out_4_2),
	.datab(lpp_ram_data_out_4_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][4]~22_combout ),
	.cout());
defparam \ram_in_reg[6][4]~22 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][4]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][4]~23 (
	.dataa(lpp_ram_data_out_4_0),
	.datab(lpp_ram_data_out_4_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][4]~23_combout ),
	.cout());
defparam \ram_in_reg[4][4]~23 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][4]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][3]~14 (
	.dataa(lpp_ram_data_out_3_2),
	.datab(lpp_ram_data_out_3_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][3]~14_combout ),
	.cout());
defparam \ram_in_reg[6][3]~14 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][3]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][3]~15 (
	.dataa(lpp_ram_data_out_3_0),
	.datab(lpp_ram_data_out_3_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][3]~15_combout ),
	.cout());
defparam \ram_in_reg[4][3]~15 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][3]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][2]~4 (
	.dataa(lpp_ram_data_out_12_2),
	.datab(lpp_ram_data_out_12_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][2]~4_combout ),
	.cout());
defparam \ram_in_reg[2][2]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][2]~5 (
	.dataa(lpp_ram_data_out_12_0),
	.datab(lpp_ram_data_out_12_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][2]~5_combout ),
	.cout());
defparam \ram_in_reg[0][2]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][1]~68 (
	.dataa(lpp_ram_data_out_11_2),
	.datab(lpp_ram_data_out_11_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~68_combout ),
	.cout());
defparam \ram_in_reg[2][1]~68 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][1]~69 (
	.dataa(lpp_ram_data_out_11_0),
	.datab(lpp_ram_data_out_11_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~69_combout ),
	.cout());
defparam \ram_in_reg[0][1]~69 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][0]~76 (
	.dataa(lpp_ram_data_out_10_2),
	.datab(lpp_ram_data_out_10_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][0]~76_combout ),
	.cout());
defparam \ram_in_reg[2][0]~76 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][0]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][0]~77 (
	.dataa(lpp_ram_data_out_10_0),
	.datab(lpp_ram_data_out_10_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][0]~77_combout ),
	.cout());
defparam \ram_in_reg[0][0]~77 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][0]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][9]~60 (
	.dataa(lpp_ram_data_out_19_2),
	.datab(lpp_ram_data_out_19_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][9]~60_combout ),
	.cout());
defparam \ram_in_reg[2][9]~60 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][9]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][9]~61 (
	.dataa(lpp_ram_data_out_19_0),
	.datab(lpp_ram_data_out_19_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][9]~61_combout ),
	.cout());
defparam \ram_in_reg[0][9]~61 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][9]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][8]~52 (
	.dataa(lpp_ram_data_out_18_2),
	.datab(lpp_ram_data_out_18_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][8]~52_combout ),
	.cout());
defparam \ram_in_reg[2][8]~52 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][8]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][8]~53 (
	.dataa(lpp_ram_data_out_18_0),
	.datab(lpp_ram_data_out_18_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][8]~53_combout ),
	.cout());
defparam \ram_in_reg[0][8]~53 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][8]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][7]~44 (
	.dataa(lpp_ram_data_out_17_2),
	.datab(lpp_ram_data_out_17_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][7]~44_combout ),
	.cout());
defparam \ram_in_reg[2][7]~44 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][7]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][7]~45 (
	.dataa(lpp_ram_data_out_17_0),
	.datab(lpp_ram_data_out_17_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][7]~45_combout ),
	.cout());
defparam \ram_in_reg[0][7]~45 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][7]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][6]~36 (
	.dataa(lpp_ram_data_out_16_2),
	.datab(lpp_ram_data_out_16_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][6]~36_combout ),
	.cout());
defparam \ram_in_reg[2][6]~36 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][6]~37 (
	.dataa(lpp_ram_data_out_16_0),
	.datab(lpp_ram_data_out_16_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][6]~37_combout ),
	.cout());
defparam \ram_in_reg[0][6]~37 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][6]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][5]~28 (
	.dataa(lpp_ram_data_out_15_2),
	.datab(lpp_ram_data_out_15_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~28_combout ),
	.cout());
defparam \ram_in_reg[2][5]~28 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][5]~29 (
	.dataa(lpp_ram_data_out_15_0),
	.datab(lpp_ram_data_out_15_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~29_combout ),
	.cout());
defparam \ram_in_reg[0][5]~29 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][4]~20 (
	.dataa(lpp_ram_data_out_14_2),
	.datab(lpp_ram_data_out_14_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][4]~20_combout ),
	.cout());
defparam \ram_in_reg[2][4]~20 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][4]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][4]~21 (
	.dataa(lpp_ram_data_out_14_0),
	.datab(lpp_ram_data_out_14_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][4]~21_combout ),
	.cout());
defparam \ram_in_reg[0][4]~21 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][4]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][3]~12 (
	.dataa(lpp_ram_data_out_13_2),
	.datab(lpp_ram_data_out_13_3),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~12_combout ),
	.cout());
defparam \ram_in_reg[2][3]~12 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][3]~13 (
	.dataa(lpp_ram_data_out_13_0),
	.datab(lpp_ram_data_out_13_1),
	.datac(gnd),
	.datad(tdl_arr_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~13_combout ),
	.cout());
defparam \ram_in_reg[0][3]~13 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~13 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cxb_data_r_1 (
	ram_in_reg_7_0,
	ram_in_reg_5_0,
	ram_in_reg_6_0,
	ram_in_reg_8_0,
	ram_in_reg_4_0,
	ram_in_reg_7_2,
	ram_in_reg_5_2,
	ram_in_reg_6_2,
	ram_in_reg_8_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_3_0,
	ram_in_reg_2_2,
	ram_in_reg_2_0,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	ram_in_reg_0_2,
	ram_in_reg_0_0,
	ram_in_reg_7_1,
	ram_in_reg_5_1,
	ram_in_reg_6_1,
	ram_in_reg_8_1,
	ram_in_reg_4_1,
	ram_in_reg_7_3,
	ram_in_reg_5_3,
	ram_in_reg_6_3,
	ram_in_reg_8_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_3_1,
	ram_in_reg_2_3,
	ram_in_reg_2_1,
	ram_in_reg_1_3,
	ram_in_reg_1_1,
	ram_in_reg_0_3,
	ram_in_reg_0_1,
	ram_in_reg_9_0,
	ram_in_reg_9_2,
	ram_in_reg_9_1,
	ram_in_reg_9_3,
	ram_in_reg_5_4,
	ram_in_reg_6_4,
	ram_in_reg_7_4,
	ram_in_reg_8_4,
	ram_in_reg_4_4,
	ram_in_reg_5_6,
	ram_in_reg_6_6,
	ram_in_reg_7_6,
	ram_in_reg_8_6,
	ram_in_reg_4_6,
	ram_in_reg_3_6,
	ram_in_reg_3_4,
	ram_in_reg_2_6,
	ram_in_reg_2_4,
	ram_in_reg_1_6,
	ram_in_reg_1_4,
	ram_in_reg_0_6,
	ram_in_reg_0_4,
	ram_in_reg_5_5,
	ram_in_reg_6_5,
	ram_in_reg_7_5,
	ram_in_reg_8_5,
	ram_in_reg_4_5,
	ram_in_reg_5_7,
	ram_in_reg_6_7,
	ram_in_reg_7_7,
	ram_in_reg_8_7,
	ram_in_reg_4_7,
	ram_in_reg_3_7,
	ram_in_reg_3_5,
	ram_in_reg_2_7,
	ram_in_reg_2_5,
	ram_in_reg_1_7,
	ram_in_reg_1_5,
	ram_in_reg_0_7,
	ram_in_reg_0_5,
	ram_in_reg_9_4,
	ram_in_reg_9_6,
	ram_in_reg_9_5,
	ram_in_reg_9_7,
	global_clock_enable,
	ram_data_out0_17,
	ram_data_out1_17,
	sw_r_tdl_0_4,
	ram_data_out2_17,
	ram_data_out3_17,
	sw_r_tdl_1_4,
	ram_data_out0_15,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_16,
	ram_data_out1_16,
	ram_data_out2_16,
	ram_data_out3_16,
	ram_data_out0_18,
	ram_data_out1_18,
	ram_data_out2_18,
	ram_data_out3_18,
	ram_data_out0_14,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_13,
	ram_data_out1_13,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_12,
	ram_data_out1_12,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_11,
	ram_data_out1_11,
	ram_data_out2_10,
	ram_data_out3_10,
	ram_data_out0_10,
	ram_data_out1_10,
	ram_data_out0_19,
	ram_data_out1_19,
	ram_data_out2_19,
	ram_data_out3_19,
	ram_data_out0_5,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_6,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_7,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_4,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_3,
	ram_data_out1_3,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_2,
	ram_data_out1_2,
	ram_data_out2_1,
	ram_data_out3_1,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_0,
	ram_data_out3_0,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out2_9,
	ram_data_out3_9,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_in_reg_7_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_6_0;
output 	ram_in_reg_8_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_7_2;
output 	ram_in_reg_5_2;
output 	ram_in_reg_6_2;
output 	ram_in_reg_8_2;
output 	ram_in_reg_4_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_0;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_0;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_0;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_0;
output 	ram_in_reg_7_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_6_1;
output 	ram_in_reg_8_1;
output 	ram_in_reg_4_1;
output 	ram_in_reg_7_3;
output 	ram_in_reg_5_3;
output 	ram_in_reg_6_3;
output 	ram_in_reg_8_3;
output 	ram_in_reg_4_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_1;
output 	ram_in_reg_2_3;
output 	ram_in_reg_2_1;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_1;
output 	ram_in_reg_0_3;
output 	ram_in_reg_0_1;
output 	ram_in_reg_9_0;
output 	ram_in_reg_9_2;
output 	ram_in_reg_9_1;
output 	ram_in_reg_9_3;
output 	ram_in_reg_5_4;
output 	ram_in_reg_6_4;
output 	ram_in_reg_7_4;
output 	ram_in_reg_8_4;
output 	ram_in_reg_4_4;
output 	ram_in_reg_5_6;
output 	ram_in_reg_6_6;
output 	ram_in_reg_7_6;
output 	ram_in_reg_8_6;
output 	ram_in_reg_4_6;
output 	ram_in_reg_3_6;
output 	ram_in_reg_3_4;
output 	ram_in_reg_2_6;
output 	ram_in_reg_2_4;
output 	ram_in_reg_1_6;
output 	ram_in_reg_1_4;
output 	ram_in_reg_0_6;
output 	ram_in_reg_0_4;
output 	ram_in_reg_5_5;
output 	ram_in_reg_6_5;
output 	ram_in_reg_7_5;
output 	ram_in_reg_8_5;
output 	ram_in_reg_4_5;
output 	ram_in_reg_5_7;
output 	ram_in_reg_6_7;
output 	ram_in_reg_7_7;
output 	ram_in_reg_8_7;
output 	ram_in_reg_4_7;
output 	ram_in_reg_3_7;
output 	ram_in_reg_3_5;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_5;
output 	ram_in_reg_1_7;
output 	ram_in_reg_1_5;
output 	ram_in_reg_0_7;
output 	ram_in_reg_0_5;
output 	ram_in_reg_9_4;
output 	ram_in_reg_9_6;
output 	ram_in_reg_9_5;
output 	ram_in_reg_9_7;
input 	global_clock_enable;
input 	ram_data_out0_17;
input 	ram_data_out1_17;
input 	sw_r_tdl_0_4;
input 	ram_data_out2_17;
input 	ram_data_out3_17;
input 	sw_r_tdl_1_4;
input 	ram_data_out0_15;
input 	ram_data_out1_15;
input 	ram_data_out2_15;
input 	ram_data_out3_15;
input 	ram_data_out0_16;
input 	ram_data_out1_16;
input 	ram_data_out2_16;
input 	ram_data_out3_16;
input 	ram_data_out0_18;
input 	ram_data_out1_18;
input 	ram_data_out2_18;
input 	ram_data_out3_18;
input 	ram_data_out0_14;
input 	ram_data_out1_14;
input 	ram_data_out2_14;
input 	ram_data_out3_14;
input 	ram_data_out2_13;
input 	ram_data_out3_13;
input 	ram_data_out0_13;
input 	ram_data_out1_13;
input 	ram_data_out2_12;
input 	ram_data_out3_12;
input 	ram_data_out0_12;
input 	ram_data_out1_12;
input 	ram_data_out2_11;
input 	ram_data_out3_11;
input 	ram_data_out0_11;
input 	ram_data_out1_11;
input 	ram_data_out2_10;
input 	ram_data_out3_10;
input 	ram_data_out0_10;
input 	ram_data_out1_10;
input 	ram_data_out0_19;
input 	ram_data_out1_19;
input 	ram_data_out2_19;
input 	ram_data_out3_19;
input 	ram_data_out0_5;
input 	ram_data_out1_5;
input 	ram_data_out2_5;
input 	ram_data_out3_5;
input 	ram_data_out0_6;
input 	ram_data_out1_6;
input 	ram_data_out2_6;
input 	ram_data_out3_6;
input 	ram_data_out0_7;
input 	ram_data_out1_7;
input 	ram_data_out2_7;
input 	ram_data_out3_7;
input 	ram_data_out0_8;
input 	ram_data_out1_8;
input 	ram_data_out2_8;
input 	ram_data_out3_8;
input 	ram_data_out0_4;
input 	ram_data_out1_4;
input 	ram_data_out2_4;
input 	ram_data_out3_4;
input 	ram_data_out2_3;
input 	ram_data_out3_3;
input 	ram_data_out0_3;
input 	ram_data_out1_3;
input 	ram_data_out2_2;
input 	ram_data_out3_2;
input 	ram_data_out0_2;
input 	ram_data_out1_2;
input 	ram_data_out2_1;
input 	ram_data_out3_1;
input 	ram_data_out0_1;
input 	ram_data_out1_1;
input 	ram_data_out2_0;
input 	ram_data_out3_0;
input 	ram_data_out0_0;
input 	ram_data_out1_0;
input 	ram_data_out0_9;
input 	ram_data_out1_9;
input 	ram_data_out2_9;
input 	ram_data_out3_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[0][7]~0_combout ;
wire \ram_in_reg[2][7]~5_combout ;
wire \ram_in_reg[0][5]~2_combout ;
wire \ram_in_reg[2][5]~7_combout ;
wire \ram_in_reg[0][6]~1_combout ;
wire \ram_in_reg[2][6]~6_combout ;
wire \ram_in_reg[0][8]~3_combout ;
wire \ram_in_reg[2][8]~8_combout ;
wire \ram_in_reg[0][4]~4_combout ;
wire \ram_in_reg[2][4]~9_combout ;
wire \ram_in_reg[2][3]~76_combout ;
wire \ram_in_reg[0][3]~77_combout ;
wire \ram_in_reg[2][2]~64_combout ;
wire \ram_in_reg[0][2]~67_combout ;
wire \ram_in_reg[2][1]~65_combout ;
wire \ram_in_reg[0][1]~68_combout ;
wire \ram_in_reg[2][0]~66_combout ;
wire \ram_in_reg[0][0]~69_combout ;
wire \ram_in_reg[1][7]~10_combout ;
wire \ram_in_reg[3][7]~15_combout ;
wire \ram_in_reg[1][5]~12_combout ;
wire \ram_in_reg[3][5]~17_combout ;
wire \ram_in_reg[1][6]~11_combout ;
wire \ram_in_reg[3][6]~16_combout ;
wire \ram_in_reg[1][8]~13_combout ;
wire \ram_in_reg[3][8]~18_combout ;
wire \ram_in_reg[1][4]~14_combout ;
wire \ram_in_reg[3][4]~19_combout ;
wire \ram_in_reg[3][3]~62_combout ;
wire \ram_in_reg[1][3]~63_combout ;
wire \ram_in_reg[3][2]~54_combout ;
wire \ram_in_reg[1][2]~57_combout ;
wire \ram_in_reg[3][1]~55_combout ;
wire \ram_in_reg[1][1]~58_combout ;
wire \ram_in_reg[3][0]~56_combout ;
wire \ram_in_reg[1][0]~59_combout ;
wire \ram_in_reg[0][9]~20_combout ;
wire \ram_in_reg[2][9]~21_combout ;
wire \ram_in_reg[1][9]~22_combout ;
wire \ram_in_reg[3][9]~23_combout ;
wire \ram_in_reg[4][5]~25_combout ;
wire \ram_in_reg[6][5]~30_combout ;
wire \ram_in_reg[4][6]~24_combout ;
wire \ram_in_reg[6][6]~29_combout ;
wire \ram_in_reg[4][7]~26_combout ;
wire \ram_in_reg[6][7]~31_combout ;
wire \ram_in_reg[4][8]~27_combout ;
wire \ram_in_reg[6][8]~32_combout ;
wire \ram_in_reg[4][4]~28_combout ;
wire \ram_in_reg[6][4]~33_combout ;
wire \ram_in_reg[6][3]~60_combout ;
wire \ram_in_reg[4][3]~61_combout ;
wire \ram_in_reg[6][2]~48_combout ;
wire \ram_in_reg[4][2]~51_combout ;
wire \ram_in_reg[6][1]~49_combout ;
wire \ram_in_reg[4][1]~52_combout ;
wire \ram_in_reg[6][0]~50_combout ;
wire \ram_in_reg[4][0]~53_combout ;
wire \ram_in_reg[5][5]~35_combout ;
wire \ram_in_reg[7][5]~40_combout ;
wire \ram_in_reg[5][6]~34_combout ;
wire \ram_in_reg[7][6]~39_combout ;
wire \ram_in_reg[5][7]~36_combout ;
wire \ram_in_reg[7][7]~41_combout ;
wire \ram_in_reg[5][8]~37_combout ;
wire \ram_in_reg[7][8]~42_combout ;
wire \ram_in_reg[5][4]~38_combout ;
wire \ram_in_reg[7][4]~43_combout ;
wire \ram_in_reg[7][3]~78_combout ;
wire \ram_in_reg[5][3]~79_combout ;
wire \ram_in_reg[7][2]~70_combout ;
wire \ram_in_reg[5][2]~73_combout ;
wire \ram_in_reg[7][1]~71_combout ;
wire \ram_in_reg[5][1]~74_combout ;
wire \ram_in_reg[7][0]~72_combout ;
wire \ram_in_reg[5][0]~75_combout ;
wire \ram_in_reg[4][9]~44_combout ;
wire \ram_in_reg[6][9]~45_combout ;
wire \ram_in_reg[5][9]~46_combout ;
wire \ram_in_reg[7][9]~47_combout ;


dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\ram_in_reg[0][7]~0_combout ),
	.asdata(\ram_in_reg[2][7]~5_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\ram_in_reg[0][5]~2_combout ),
	.asdata(\ram_in_reg[2][5]~7_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\ram_in_reg[0][6]~1_combout ),
	.asdata(\ram_in_reg[2][6]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[0][8] (
	.clk(clk),
	.d(\ram_in_reg[0][8]~3_combout ),
	.asdata(\ram_in_reg[2][8]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_0),
	.prn(vcc));
defparam \ram_in_reg[0][8] .is_wysiwyg = "true";
defparam \ram_in_reg[0][8] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\ram_in_reg[0][4]~4_combout ),
	.asdata(\ram_in_reg[2][4]~9_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\ram_in_reg[2][7]~5_combout ),
	.asdata(\ram_in_reg[0][7]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\ram_in_reg[2][5]~7_combout ),
	.asdata(\ram_in_reg[0][5]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\ram_in_reg[2][6]~6_combout ),
	.asdata(\ram_in_reg[0][6]~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[2][8] (
	.clk(clk),
	.d(\ram_in_reg[2][8]~8_combout ),
	.asdata(\ram_in_reg[0][8]~3_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_2),
	.prn(vcc));
defparam \ram_in_reg[2][8] .is_wysiwyg = "true";
defparam \ram_in_reg[2][8] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\ram_in_reg[2][4]~9_combout ),
	.asdata(\ram_in_reg[0][4]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\ram_in_reg[2][3]~76_combout ),
	.asdata(\ram_in_reg[0][3]~77_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\ram_in_reg[0][3]~77_combout ),
	.asdata(\ram_in_reg[2][3]~76_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\ram_in_reg[2][2]~64_combout ),
	.asdata(\ram_in_reg[0][2]~67_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\ram_in_reg[0][2]~67_combout ),
	.asdata(\ram_in_reg[2][2]~64_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\ram_in_reg[2][1]~65_combout ),
	.asdata(\ram_in_reg[0][1]~68_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\ram_in_reg[0][1]~68_combout ),
	.asdata(\ram_in_reg[2][1]~65_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\ram_in_reg[2][0]~66_combout ),
	.asdata(\ram_in_reg[0][0]~69_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\ram_in_reg[0][0]~69_combout ),
	.asdata(\ram_in_reg[2][0]~66_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\ram_in_reg[1][7]~10_combout ),
	.asdata(\ram_in_reg[3][7]~15_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\ram_in_reg[1][5]~12_combout ),
	.asdata(\ram_in_reg[3][5]~17_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\ram_in_reg[1][6]~11_combout ),
	.asdata(\ram_in_reg[3][6]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[1][8] (
	.clk(clk),
	.d(\ram_in_reg[1][8]~13_combout ),
	.asdata(\ram_in_reg[3][8]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_1),
	.prn(vcc));
defparam \ram_in_reg[1][8] .is_wysiwyg = "true";
defparam \ram_in_reg[1][8] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\ram_in_reg[1][4]~14_combout ),
	.asdata(\ram_in_reg[3][4]~19_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\ram_in_reg[3][7]~15_combout ),
	.asdata(\ram_in_reg[1][7]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\ram_in_reg[3][5]~17_combout ),
	.asdata(\ram_in_reg[1][5]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\ram_in_reg[3][6]~16_combout ),
	.asdata(\ram_in_reg[1][6]~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[3][8] (
	.clk(clk),
	.d(\ram_in_reg[3][8]~18_combout ),
	.asdata(\ram_in_reg[1][8]~13_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_3),
	.prn(vcc));
defparam \ram_in_reg[3][8] .is_wysiwyg = "true";
defparam \ram_in_reg[3][8] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\ram_in_reg[3][4]~19_combout ),
	.asdata(\ram_in_reg[1][4]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~62_combout ),
	.asdata(\ram_in_reg[1][3]~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\ram_in_reg[1][3]~63_combout ),
	.asdata(\ram_in_reg[3][3]~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\ram_in_reg[3][2]~54_combout ),
	.asdata(\ram_in_reg[1][2]~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~57_combout ),
	.asdata(\ram_in_reg[3][2]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\ram_in_reg[3][1]~55_combout ),
	.asdata(\ram_in_reg[1][1]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\ram_in_reg[1][1]~58_combout ),
	.asdata(\ram_in_reg[3][1]~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\ram_in_reg[3][0]~56_combout ),
	.asdata(\ram_in_reg[1][0]~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\ram_in_reg[1][0]~59_combout ),
	.asdata(\ram_in_reg[3][0]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[0][9] (
	.clk(clk),
	.d(\ram_in_reg[0][9]~20_combout ),
	.asdata(\ram_in_reg[2][9]~21_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_0),
	.prn(vcc));
defparam \ram_in_reg[0][9] .is_wysiwyg = "true";
defparam \ram_in_reg[0][9] .power_up = "low";

dffeas \ram_in_reg[2][9] (
	.clk(clk),
	.d(\ram_in_reg[2][9]~21_combout ),
	.asdata(\ram_in_reg[0][9]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_2),
	.prn(vcc));
defparam \ram_in_reg[2][9] .is_wysiwyg = "true";
defparam \ram_in_reg[2][9] .power_up = "low";

dffeas \ram_in_reg[1][9] (
	.clk(clk),
	.d(\ram_in_reg[1][9]~22_combout ),
	.asdata(\ram_in_reg[3][9]~23_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_1),
	.prn(vcc));
defparam \ram_in_reg[1][9] .is_wysiwyg = "true";
defparam \ram_in_reg[1][9] .power_up = "low";

dffeas \ram_in_reg[3][9] (
	.clk(clk),
	.d(\ram_in_reg[3][9]~23_combout ),
	.asdata(\ram_in_reg[1][9]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_3),
	.prn(vcc));
defparam \ram_in_reg[3][9] .is_wysiwyg = "true";
defparam \ram_in_reg[3][9] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\ram_in_reg[4][5]~25_combout ),
	.asdata(\ram_in_reg[6][5]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\ram_in_reg[4][6]~24_combout ),
	.asdata(\ram_in_reg[6][6]~29_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\ram_in_reg[4][7]~26_combout ),
	.asdata(\ram_in_reg[6][7]~31_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[4][8] (
	.clk(clk),
	.d(\ram_in_reg[4][8]~27_combout ),
	.asdata(\ram_in_reg[6][8]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_4),
	.prn(vcc));
defparam \ram_in_reg[4][8] .is_wysiwyg = "true";
defparam \ram_in_reg[4][8] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\ram_in_reg[4][4]~28_combout ),
	.asdata(\ram_in_reg[6][4]~33_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\ram_in_reg[6][5]~30_combout ),
	.asdata(\ram_in_reg[4][5]~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\ram_in_reg[6][6]~29_combout ),
	.asdata(\ram_in_reg[4][6]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\ram_in_reg[6][7]~31_combout ),
	.asdata(\ram_in_reg[4][7]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[6][8] (
	.clk(clk),
	.d(\ram_in_reg[6][8]~32_combout ),
	.asdata(\ram_in_reg[4][8]~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_6),
	.prn(vcc));
defparam \ram_in_reg[6][8] .is_wysiwyg = "true";
defparam \ram_in_reg[6][8] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\ram_in_reg[6][4]~33_combout ),
	.asdata(\ram_in_reg[4][4]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\ram_in_reg[6][3]~60_combout ),
	.asdata(\ram_in_reg[4][3]~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\ram_in_reg[4][3]~61_combout ),
	.asdata(\ram_in_reg[6][3]~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\ram_in_reg[6][2]~48_combout ),
	.asdata(\ram_in_reg[4][2]~51_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\ram_in_reg[4][2]~51_combout ),
	.asdata(\ram_in_reg[6][2]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\ram_in_reg[6][1]~49_combout ),
	.asdata(\ram_in_reg[4][1]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\ram_in_reg[4][1]~52_combout ),
	.asdata(\ram_in_reg[6][1]~49_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\ram_in_reg[6][0]~50_combout ),
	.asdata(\ram_in_reg[4][0]~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\ram_in_reg[4][0]~53_combout ),
	.asdata(\ram_in_reg[6][0]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\ram_in_reg[5][5]~35_combout ),
	.asdata(\ram_in_reg[7][5]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\ram_in_reg[5][6]~34_combout ),
	.asdata(\ram_in_reg[7][6]~39_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\ram_in_reg[5][7]~36_combout ),
	.asdata(\ram_in_reg[7][7]~41_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[5][8] (
	.clk(clk),
	.d(\ram_in_reg[5][8]~37_combout ),
	.asdata(\ram_in_reg[7][8]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_5),
	.prn(vcc));
defparam \ram_in_reg[5][8] .is_wysiwyg = "true";
defparam \ram_in_reg[5][8] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\ram_in_reg[5][4]~38_combout ),
	.asdata(\ram_in_reg[7][4]~43_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\ram_in_reg[7][5]~40_combout ),
	.asdata(\ram_in_reg[5][5]~35_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\ram_in_reg[7][6]~39_combout ),
	.asdata(\ram_in_reg[5][6]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\ram_in_reg[7][7]~41_combout ),
	.asdata(\ram_in_reg[5][7]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[7][8] (
	.clk(clk),
	.d(\ram_in_reg[7][8]~42_combout ),
	.asdata(\ram_in_reg[5][8]~37_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_8_7),
	.prn(vcc));
defparam \ram_in_reg[7][8] .is_wysiwyg = "true";
defparam \ram_in_reg[7][8] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\ram_in_reg[7][4]~43_combout ),
	.asdata(\ram_in_reg[5][4]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\ram_in_reg[7][3]~78_combout ),
	.asdata(\ram_in_reg[5][3]~79_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\ram_in_reg[5][3]~79_combout ),
	.asdata(\ram_in_reg[7][3]~78_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\ram_in_reg[7][2]~70_combout ),
	.asdata(\ram_in_reg[5][2]~73_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\ram_in_reg[5][2]~73_combout ),
	.asdata(\ram_in_reg[7][2]~70_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\ram_in_reg[7][1]~71_combout ),
	.asdata(\ram_in_reg[5][1]~74_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\ram_in_reg[5][1]~74_combout ),
	.asdata(\ram_in_reg[7][1]~71_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\ram_in_reg[7][0]~72_combout ),
	.asdata(\ram_in_reg[5][0]~75_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\ram_in_reg[5][0]~75_combout ),
	.asdata(\ram_in_reg[7][0]~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[4][9] (
	.clk(clk),
	.d(\ram_in_reg[4][9]~44_combout ),
	.asdata(\ram_in_reg[6][9]~45_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_4),
	.prn(vcc));
defparam \ram_in_reg[4][9] .is_wysiwyg = "true";
defparam \ram_in_reg[4][9] .power_up = "low";

dffeas \ram_in_reg[6][9] (
	.clk(clk),
	.d(\ram_in_reg[6][9]~45_combout ),
	.asdata(\ram_in_reg[4][9]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_6),
	.prn(vcc));
defparam \ram_in_reg[6][9] .is_wysiwyg = "true";
defparam \ram_in_reg[6][9] .power_up = "low";

dffeas \ram_in_reg[5][9] (
	.clk(clk),
	.d(\ram_in_reg[5][9]~46_combout ),
	.asdata(\ram_in_reg[7][9]~47_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_5),
	.prn(vcc));
defparam \ram_in_reg[5][9] .is_wysiwyg = "true";
defparam \ram_in_reg[5][9] .power_up = "low";

dffeas \ram_in_reg[7][9] (
	.clk(clk),
	.d(\ram_in_reg[7][9]~47_combout ),
	.asdata(\ram_in_reg[5][9]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(sw_r_tdl_1_4),
	.ena(global_clock_enable),
	.q(ram_in_reg_9_7),
	.prn(vcc));
defparam \ram_in_reg[7][9] .is_wysiwyg = "true";
defparam \ram_in_reg[7][9] .power_up = "low";

cycloneive_lcell_comb \ram_in_reg[0][7]~0 (
	.dataa(ram_data_out0_17),
	.datab(ram_data_out1_17),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][7]~0_combout ),
	.cout());
defparam \ram_in_reg[0][7]~0 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][7]~5 (
	.dataa(ram_data_out2_17),
	.datab(ram_data_out3_17),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][7]~5_combout ),
	.cout());
defparam \ram_in_reg[2][7]~5 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][7]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][5]~2 (
	.dataa(ram_data_out0_15),
	.datab(ram_data_out1_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][5]~2_combout ),
	.cout());
defparam \ram_in_reg[0][5]~2 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][5]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][5]~7 (
	.dataa(ram_data_out2_15),
	.datab(ram_data_out3_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][5]~7_combout ),
	.cout());
defparam \ram_in_reg[2][5]~7 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][5]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][6]~1 (
	.dataa(ram_data_out0_16),
	.datab(ram_data_out1_16),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][6]~1_combout ),
	.cout());
defparam \ram_in_reg[0][6]~1 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][6]~6 (
	.dataa(ram_data_out2_16),
	.datab(ram_data_out3_16),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][6]~6_combout ),
	.cout());
defparam \ram_in_reg[2][6]~6 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][8]~3 (
	.dataa(ram_data_out0_18),
	.datab(ram_data_out1_18),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][8]~3_combout ),
	.cout());
defparam \ram_in_reg[0][8]~3 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][8]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][8]~8 (
	.dataa(ram_data_out2_18),
	.datab(ram_data_out3_18),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][8]~8_combout ),
	.cout());
defparam \ram_in_reg[2][8]~8 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][8]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][4]~4 (
	.dataa(ram_data_out0_14),
	.datab(ram_data_out1_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][4]~4_combout ),
	.cout());
defparam \ram_in_reg[0][4]~4 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][4]~9 (
	.dataa(ram_data_out2_14),
	.datab(ram_data_out3_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][4]~9_combout ),
	.cout());
defparam \ram_in_reg[2][4]~9 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][4]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][3]~76 (
	.dataa(ram_data_out2_13),
	.datab(ram_data_out3_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][3]~76_combout ),
	.cout());
defparam \ram_in_reg[2][3]~76 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][3]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][3]~77 (
	.dataa(ram_data_out0_13),
	.datab(ram_data_out1_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][3]~77_combout ),
	.cout());
defparam \ram_in_reg[0][3]~77 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][3]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][2]~64 (
	.dataa(ram_data_out2_12),
	.datab(ram_data_out3_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][2]~64_combout ),
	.cout());
defparam \ram_in_reg[2][2]~64 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][2]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][2]~67 (
	.dataa(ram_data_out0_12),
	.datab(ram_data_out1_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][2]~67_combout ),
	.cout());
defparam \ram_in_reg[0][2]~67 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][2]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][1]~65 (
	.dataa(ram_data_out2_11),
	.datab(ram_data_out3_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][1]~65_combout ),
	.cout());
defparam \ram_in_reg[2][1]~65 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][1]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][1]~68 (
	.dataa(ram_data_out0_11),
	.datab(ram_data_out1_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][1]~68_combout ),
	.cout());
defparam \ram_in_reg[0][1]~68 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][1]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][0]~66 (
	.dataa(ram_data_out2_10),
	.datab(ram_data_out3_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][0]~66_combout ),
	.cout());
defparam \ram_in_reg[2][0]~66 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][0]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][0]~69 (
	.dataa(ram_data_out0_10),
	.datab(ram_data_out1_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][0]~69_combout ),
	.cout());
defparam \ram_in_reg[0][0]~69 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][0]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][7]~10 (
	.dataa(ram_data_out1_17),
	.datab(ram_data_out2_17),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][7]~10_combout ),
	.cout());
defparam \ram_in_reg[1][7]~10 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][7]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][7]~15 (
	.dataa(ram_data_out3_17),
	.datab(ram_data_out0_17),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][7]~15_combout ),
	.cout());
defparam \ram_in_reg[3][7]~15 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][5]~12 (
	.dataa(ram_data_out1_15),
	.datab(ram_data_out2_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][5]~12_combout ),
	.cout());
defparam \ram_in_reg[1][5]~12 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][5]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][5]~17 (
	.dataa(ram_data_out3_15),
	.datab(ram_data_out0_15),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][5]~17_combout ),
	.cout());
defparam \ram_in_reg[3][5]~17 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][5]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][6]~11 (
	.dataa(ram_data_out1_16),
	.datab(ram_data_out2_16),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][6]~11_combout ),
	.cout());
defparam \ram_in_reg[1][6]~11 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][6]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][6]~16 (
	.dataa(ram_data_out3_16),
	.datab(ram_data_out0_16),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][6]~16_combout ),
	.cout());
defparam \ram_in_reg[3][6]~16 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][6]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][8]~13 (
	.dataa(ram_data_out1_18),
	.datab(ram_data_out2_18),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][8]~13_combout ),
	.cout());
defparam \ram_in_reg[1][8]~13 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][8]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][8]~18 (
	.dataa(ram_data_out3_18),
	.datab(ram_data_out0_18),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][8]~18_combout ),
	.cout());
defparam \ram_in_reg[3][8]~18 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][8]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][4]~14 (
	.dataa(ram_data_out1_14),
	.datab(ram_data_out2_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][4]~14_combout ),
	.cout());
defparam \ram_in_reg[1][4]~14 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][4]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][4]~19 (
	.dataa(ram_data_out3_14),
	.datab(ram_data_out0_14),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][4]~19_combout ),
	.cout());
defparam \ram_in_reg[3][4]~19 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][4]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][3]~62 (
	.dataa(ram_data_out3_13),
	.datab(ram_data_out0_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][3]~62_combout ),
	.cout());
defparam \ram_in_reg[3][3]~62 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][3]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][3]~63 (
	.dataa(ram_data_out1_13),
	.datab(ram_data_out2_13),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][3]~63_combout ),
	.cout());
defparam \ram_in_reg[1][3]~63 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][3]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][2]~54 (
	.dataa(ram_data_out3_12),
	.datab(ram_data_out0_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][2]~54_combout ),
	.cout());
defparam \ram_in_reg[3][2]~54 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][2]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][2]~57 (
	.dataa(ram_data_out1_12),
	.datab(ram_data_out2_12),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][2]~57_combout ),
	.cout());
defparam \ram_in_reg[1][2]~57 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][2]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][1]~55 (
	.dataa(ram_data_out3_11),
	.datab(ram_data_out0_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][1]~55_combout ),
	.cout());
defparam \ram_in_reg[3][1]~55 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][1]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][1]~58 (
	.dataa(ram_data_out1_11),
	.datab(ram_data_out2_11),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][1]~58_combout ),
	.cout());
defparam \ram_in_reg[1][1]~58 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][1]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][0]~56 (
	.dataa(ram_data_out3_10),
	.datab(ram_data_out0_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][0]~56_combout ),
	.cout());
defparam \ram_in_reg[3][0]~56 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][0]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][0]~59 (
	.dataa(ram_data_out1_10),
	.datab(ram_data_out2_10),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][0]~59_combout ),
	.cout());
defparam \ram_in_reg[1][0]~59 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][0]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[0][9]~20 (
	.dataa(ram_data_out0_19),
	.datab(ram_data_out1_19),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[0][9]~20_combout ),
	.cout());
defparam \ram_in_reg[0][9]~20 .lut_mask = 16'hAACC;
defparam \ram_in_reg[0][9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[2][9]~21 (
	.dataa(ram_data_out2_19),
	.datab(ram_data_out3_19),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[2][9]~21_combout ),
	.cout());
defparam \ram_in_reg[2][9]~21 .lut_mask = 16'hAACC;
defparam \ram_in_reg[2][9]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[1][9]~22 (
	.dataa(ram_data_out1_19),
	.datab(ram_data_out2_19),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[1][9]~22_combout ),
	.cout());
defparam \ram_in_reg[1][9]~22 .lut_mask = 16'hAACC;
defparam \ram_in_reg[1][9]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[3][9]~23 (
	.dataa(ram_data_out3_19),
	.datab(ram_data_out0_19),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[3][9]~23_combout ),
	.cout());
defparam \ram_in_reg[3][9]~23 .lut_mask = 16'hAACC;
defparam \ram_in_reg[3][9]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][5]~25 (
	.dataa(ram_data_out0_5),
	.datab(ram_data_out1_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][5]~25_combout ),
	.cout());
defparam \ram_in_reg[4][5]~25 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][5]~30 (
	.dataa(ram_data_out2_5),
	.datab(ram_data_out3_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][5]~30_combout ),
	.cout());
defparam \ram_in_reg[6][5]~30 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][5]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][6]~24 (
	.dataa(ram_data_out0_6),
	.datab(ram_data_out1_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][6]~24_combout ),
	.cout());
defparam \ram_in_reg[4][6]~24 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][6]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][6]~29 (
	.dataa(ram_data_out2_6),
	.datab(ram_data_out3_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][6]~29_combout ),
	.cout());
defparam \ram_in_reg[6][6]~29 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][6]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][7]~26 (
	.dataa(ram_data_out0_7),
	.datab(ram_data_out1_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][7]~26_combout ),
	.cout());
defparam \ram_in_reg[4][7]~26 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][7]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][7]~31 (
	.dataa(ram_data_out2_7),
	.datab(ram_data_out3_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][7]~31_combout ),
	.cout());
defparam \ram_in_reg[6][7]~31 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][7]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][8]~27 (
	.dataa(ram_data_out0_8),
	.datab(ram_data_out1_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][8]~27_combout ),
	.cout());
defparam \ram_in_reg[4][8]~27 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][8]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][8]~32 (
	.dataa(ram_data_out2_8),
	.datab(ram_data_out3_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][8]~32_combout ),
	.cout());
defparam \ram_in_reg[6][8]~32 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][8]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][4]~28 (
	.dataa(ram_data_out0_4),
	.datab(ram_data_out1_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][4]~28_combout ),
	.cout());
defparam \ram_in_reg[4][4]~28 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][4]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][4]~33 (
	.dataa(ram_data_out2_4),
	.datab(ram_data_out3_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][4]~33_combout ),
	.cout());
defparam \ram_in_reg[6][4]~33 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][4]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][3]~60 (
	.dataa(ram_data_out2_3),
	.datab(ram_data_out3_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][3]~60_combout ),
	.cout());
defparam \ram_in_reg[6][3]~60 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][3]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][3]~61 (
	.dataa(ram_data_out0_3),
	.datab(ram_data_out1_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][3]~61_combout ),
	.cout());
defparam \ram_in_reg[4][3]~61 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][3]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][2]~48 (
	.dataa(ram_data_out2_2),
	.datab(ram_data_out3_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][2]~48_combout ),
	.cout());
defparam \ram_in_reg[6][2]~48 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][2]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][2]~51 (
	.dataa(ram_data_out0_2),
	.datab(ram_data_out1_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][2]~51_combout ),
	.cout());
defparam \ram_in_reg[4][2]~51 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][2]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][1]~49 (
	.dataa(ram_data_out2_1),
	.datab(ram_data_out3_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][1]~49_combout ),
	.cout());
defparam \ram_in_reg[6][1]~49 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][1]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][1]~52 (
	.dataa(ram_data_out0_1),
	.datab(ram_data_out1_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][1]~52_combout ),
	.cout());
defparam \ram_in_reg[4][1]~52 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][1]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][0]~50 (
	.dataa(ram_data_out2_0),
	.datab(ram_data_out3_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][0]~50_combout ),
	.cout());
defparam \ram_in_reg[6][0]~50 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][0]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][0]~53 (
	.dataa(ram_data_out0_0),
	.datab(ram_data_out1_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][0]~53_combout ),
	.cout());
defparam \ram_in_reg[4][0]~53 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][0]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][5]~35 (
	.dataa(ram_data_out1_5),
	.datab(ram_data_out2_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][5]~35_combout ),
	.cout());
defparam \ram_in_reg[5][5]~35 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][5]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][5]~40 (
	.dataa(ram_data_out3_5),
	.datab(ram_data_out0_5),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][5]~40_combout ),
	.cout());
defparam \ram_in_reg[7][5]~40 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][5]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][6]~34 (
	.dataa(ram_data_out1_6),
	.datab(ram_data_out2_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][6]~34_combout ),
	.cout());
defparam \ram_in_reg[5][6]~34 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][6]~39 (
	.dataa(ram_data_out3_6),
	.datab(ram_data_out0_6),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][6]~39_combout ),
	.cout());
defparam \ram_in_reg[7][6]~39 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][6]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][7]~36 (
	.dataa(ram_data_out1_7),
	.datab(ram_data_out2_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][7]~36_combout ),
	.cout());
defparam \ram_in_reg[5][7]~36 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][7]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][7]~41 (
	.dataa(ram_data_out3_7),
	.datab(ram_data_out0_7),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][7]~41_combout ),
	.cout());
defparam \ram_in_reg[7][7]~41 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][7]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][8]~37 (
	.dataa(ram_data_out1_8),
	.datab(ram_data_out2_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][8]~37_combout ),
	.cout());
defparam \ram_in_reg[5][8]~37 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][8]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][8]~42 (
	.dataa(ram_data_out3_8),
	.datab(ram_data_out0_8),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][8]~42_combout ),
	.cout());
defparam \ram_in_reg[7][8]~42 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][8]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][4]~38 (
	.dataa(ram_data_out1_4),
	.datab(ram_data_out2_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][4]~38_combout ),
	.cout());
defparam \ram_in_reg[5][4]~38 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][4]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][4]~43 (
	.dataa(ram_data_out3_4),
	.datab(ram_data_out0_4),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][4]~43_combout ),
	.cout());
defparam \ram_in_reg[7][4]~43 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][4]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][3]~78 (
	.dataa(ram_data_out3_3),
	.datab(ram_data_out0_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][3]~78_combout ),
	.cout());
defparam \ram_in_reg[7][3]~78 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][3]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][3]~79 (
	.dataa(ram_data_out1_3),
	.datab(ram_data_out2_3),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][3]~79_combout ),
	.cout());
defparam \ram_in_reg[5][3]~79 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][3]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][2]~70 (
	.dataa(ram_data_out3_2),
	.datab(ram_data_out0_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][2]~70_combout ),
	.cout());
defparam \ram_in_reg[7][2]~70 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][2]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][2]~73 (
	.dataa(ram_data_out1_2),
	.datab(ram_data_out2_2),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][2]~73_combout ),
	.cout());
defparam \ram_in_reg[5][2]~73 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][2]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][1]~71 (
	.dataa(ram_data_out3_1),
	.datab(ram_data_out0_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][1]~71_combout ),
	.cout());
defparam \ram_in_reg[7][1]~71 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][1]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][1]~74 (
	.dataa(ram_data_out1_1),
	.datab(ram_data_out2_1),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][1]~74_combout ),
	.cout());
defparam \ram_in_reg[5][1]~74 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][1]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][0]~72 (
	.dataa(ram_data_out3_0),
	.datab(ram_data_out0_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][0]~72_combout ),
	.cout());
defparam \ram_in_reg[7][0]~72 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][0]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][0]~75 (
	.dataa(ram_data_out1_0),
	.datab(ram_data_out2_0),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][0]~75_combout ),
	.cout());
defparam \ram_in_reg[5][0]~75 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][0]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[4][9]~44 (
	.dataa(ram_data_out0_9),
	.datab(ram_data_out1_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[4][9]~44_combout ),
	.cout());
defparam \ram_in_reg[4][9]~44 .lut_mask = 16'hAACC;
defparam \ram_in_reg[4][9]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[6][9]~45 (
	.dataa(ram_data_out2_9),
	.datab(ram_data_out3_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[6][9]~45_combout ),
	.cout());
defparam \ram_in_reg[6][9]~45 .lut_mask = 16'hAACC;
defparam \ram_in_reg[6][9]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[5][9]~46 (
	.dataa(ram_data_out1_9),
	.datab(ram_data_out2_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[5][9]~46_combout ),
	.cout());
defparam \ram_in_reg[5][9]~46 .lut_mask = 16'hAACC;
defparam \ram_in_reg[5][9]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ram_in_reg[7][9]~47 (
	.dataa(ram_data_out3_9),
	.datab(ram_data_out0_9),
	.datac(gnd),
	.datad(sw_r_tdl_0_4),
	.cin(gnd),
	.combout(\ram_in_reg[7][9]~47_combout ),
	.cout());
defparam \ram_in_reg[7][9]~47 .lut_mask = 16'hAACC;
defparam \ram_in_reg[7][9]~47 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_dataadgen (
	global_clock_enable,
	rd_addr_c_0,
	rd_addr_d_0,
	sw_0,
	rd_addr_b_1,
	rd_addr_d_1,
	sw_1,
	rd_addr_c_2,
	rd_addr_d_2,
	rd_addr_b_3,
	rd_addr_d_3,
	rd_addr_c_4,
	rd_addr_d_4,
	rd_addr_b_5,
	rd_addr_d_5,
	rd_addr_d_6,
	rd_addr_d_7,
	p_2,
	p_0,
	p_1,
	k_count_4,
	k_count_0,
	k_count_2,
	Add1,
	Mux1,
	Mux11,
	k_count_6,
	k_count_1,
	k_count_3,
	Add0,
	k_count_5,
	Add11,
	Add12,
	Mux0,
	Mux01,
	k_count_7,
	Mux02,
	Mux12,
	Mux13,
	Mux03,
	Mux04,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	rd_addr_c_0;
output 	rd_addr_d_0;
output 	sw_0;
output 	rd_addr_b_1;
output 	rd_addr_d_1;
output 	sw_1;
output 	rd_addr_c_2;
output 	rd_addr_d_2;
output 	rd_addr_b_3;
output 	rd_addr_d_3;
output 	rd_addr_c_4;
output 	rd_addr_d_4;
output 	rd_addr_b_5;
output 	rd_addr_d_5;
output 	rd_addr_d_6;
output 	rd_addr_d_7;
input 	p_2;
input 	p_0;
input 	p_1;
input 	k_count_4;
input 	k_count_0;
input 	k_count_2;
output 	Add1;
output 	Mux1;
output 	Mux11;
input 	k_count_6;
input 	k_count_1;
input 	k_count_3;
output 	Add0;
input 	k_count_5;
output 	Add11;
output 	Add12;
output 	Mux0;
output 	Mux01;
input 	k_count_7;
input 	Mux02;
output 	Mux12;
output 	Mux13;
output 	Mux03;
output 	Mux04;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux7~2_combout ;
wire \Mux10~0_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux6~0_combout ;
wire \Mux13~0_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux9~0_combout ;
wire \Mux4~0_combout ;
wire \Mux12~0_combout ;
wire \Mux3~0_combout ;
wire \Mux8~0_combout ;
wire \Mux2~0_combout ;
wire \Mux11~0_combout ;


dffeas \rd_addr_c[0] (
	.clk(clk),
	.d(\Mux7~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_0),
	.prn(vcc));
defparam \rd_addr_c[0] .is_wysiwyg = "true";
defparam \rd_addr_c[0] .power_up = "low";

dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \sw[0] (
	.clk(clk),
	.d(\Mux1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \rd_addr_b[1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_1),
	.prn(vcc));
defparam \rd_addr_b[1] .is_wysiwyg = "true";
defparam \rd_addr_b[1] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

dffeas \sw[1] (
	.clk(clk),
	.d(\Mux0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_1),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

dffeas \rd_addr_c[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_2),
	.prn(vcc));
defparam \rd_addr_c[2] .is_wysiwyg = "true";
defparam \rd_addr_c[2] .power_up = "low";

dffeas \rd_addr_d[2] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_2),
	.prn(vcc));
defparam \rd_addr_d[2] .is_wysiwyg = "true";
defparam \rd_addr_d[2] .power_up = "low";

dffeas \rd_addr_b[3] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_3),
	.prn(vcc));
defparam \rd_addr_b[3] .is_wysiwyg = "true";
defparam \rd_addr_b[3] .power_up = "low";

dffeas \rd_addr_d[3] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_3),
	.prn(vcc));
defparam \rd_addr_d[3] .is_wysiwyg = "true";
defparam \rd_addr_d[3] .power_up = "low";

dffeas \rd_addr_c[4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_c_4),
	.prn(vcc));
defparam \rd_addr_c[4] .is_wysiwyg = "true";
defparam \rd_addr_c[4] .power_up = "low";

dffeas \rd_addr_d[4] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_4),
	.prn(vcc));
defparam \rd_addr_d[4] .is_wysiwyg = "true";
defparam \rd_addr_d[4] .power_up = "low";

dffeas \rd_addr_b[5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_b_5),
	.prn(vcc));
defparam \rd_addr_b[5] .is_wysiwyg = "true";
defparam \rd_addr_b[5] .power_up = "low";

dffeas \rd_addr_d[5] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_5),
	.prn(vcc));
defparam \rd_addr_d[5] .is_wysiwyg = "true";
defparam \rd_addr_d[5] .power_up = "low";

dffeas \rd_addr_d[6] (
	.clk(clk),
	.d(k_count_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_6),
	.prn(vcc));
defparam \rd_addr_d[6] .is_wysiwyg = "true";
defparam \rd_addr_d[6] .power_up = "low";

dffeas \rd_addr_d[7] (
	.clk(clk),
	.d(k_count_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_7),
	.prn(vcc));
defparam \rd_addr_d[7] .is_wysiwyg = "true";
defparam \rd_addr_d[7] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(k_count_4),
	.datab(k_count_0),
	.datac(k_count_2),
	.datad(gnd),
	.cin(gnd),
	.combout(Add1),
	.cout());
defparam \Add1~0 .lut_mask = 16'h9696;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(gnd),
	.datab(k_count_0),
	.datac(k_count_2),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~0 .lut_mask = 16'h3CFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(k_count_0),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux11),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAAFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(k_count_0),
	.datab(k_count_2),
	.datac(k_count_1),
	.datad(k_count_3),
	.cin(gnd),
	.combout(Add0),
	.cout());
defparam \Add0~0 .lut_mask = 16'h6996;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~1 (
	.dataa(k_count_5),
	.datab(k_count_0),
	.datac(k_count_2),
	.datad(k_count_4),
	.cin(gnd),
	.combout(Add11),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(Add0),
	.datad(Add11),
	.cin(gnd),
	.combout(Add12),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(Add0),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hAAFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(k_count_1),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux01),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hAAFF;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~5 (
	.dataa(k_count_2),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux12),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hAAFF;
defparam \Mux1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~6 (
	.dataa(k_count_4),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux13),
	.cout());
defparam \Mux1~6 .lut_mask = 16'hAAFF;
defparam \Mux1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~5 (
	.dataa(k_count_3),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux03),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hAAFF;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~6 (
	.dataa(k_count_5),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(Mux04),
	.cout());
defparam \Mux0~6 .lut_mask = 16'hAAFF;
defparam \Mux0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(gnd),
	.datab(p_1),
	.datac(p_0),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'h3FCF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(p_1),
	.datab(gnd),
	.datac(gnd),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hAAFF;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~2 (
	.dataa(k_count_0),
	.datab(k_count_2),
	.datac(\Mux7~0_combout ),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hACFF;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~0 (
	.dataa(k_count_0),
	.datab(\Mux7~0_combout ),
	.datac(k_count_2),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hFFB8;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(k_count_6),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hAAFF;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~3 (
	.dataa(Add1),
	.datab(\Mux1~2_combout ),
	.datac(Mux02),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hEFFE;
defparam \Mux1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~4 (
	.dataa(Mux11),
	.datab(Mux1),
	.datac(p_1),
	.datad(\Mux1~3_combout ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'hEFFE;
defparam \Mux1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(k_count_1),
	.datab(k_count_3),
	.datac(\Mux7~0_combout ),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hACFF;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(k_count_1),
	.datab(\Mux7~0_combout ),
	.datac(k_count_3),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFFB8;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(k_count_7),
	.datab(gnd),
	.datac(gnd),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hAAFF;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(Add12),
	.datab(\Mux0~2_combout ),
	.datac(Mux02),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hEFFE;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~4 (
	.dataa(Mux01),
	.datab(Mux0),
	.datac(p_1),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hEFFE;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(p_2),
	.datab(gnd),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hA55A;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(k_count_2),
	.datab(\Mux5~0_combout ),
	.datac(k_count_4),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hB8FF;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(k_count_2),
	.datab(p_0),
	.datac(k_count_4),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFAFC;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(k_count_3),
	.datab(\Mux5~0_combout ),
	.datac(k_count_5),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hB8FF;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~0 (
	.dataa(k_count_3),
	.datab(p_0),
	.datac(k_count_5),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFAFC;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(k_count_4),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFEFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~0 (
	.dataa(k_count_4),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hEFFF;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(k_count_5),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(k_count_5),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hEFFF;
defparam \Mux11~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_dft_bfp (
	ram_in_reg_7_0,
	ram_in_reg_5_0,
	ram_in_reg_6_0,
	ram_in_reg_8_0,
	ram_in_reg_4_0,
	ram_in_reg_7_2,
	ram_in_reg_5_2,
	ram_in_reg_6_2,
	ram_in_reg_8_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_3_0,
	ram_in_reg_2_2,
	ram_in_reg_2_0,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	ram_in_reg_0_2,
	ram_in_reg_0_0,
	ram_in_reg_7_1,
	ram_in_reg_5_1,
	ram_in_reg_6_1,
	ram_in_reg_8_1,
	ram_in_reg_4_1,
	ram_in_reg_7_3,
	ram_in_reg_5_3,
	ram_in_reg_6_3,
	ram_in_reg_8_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_3_1,
	ram_in_reg_2_3,
	ram_in_reg_2_1,
	ram_in_reg_1_3,
	ram_in_reg_1_1,
	ram_in_reg_0_3,
	ram_in_reg_0_1,
	ram_in_reg_9_0,
	ram_in_reg_9_2,
	ram_in_reg_9_1,
	ram_in_reg_9_3,
	ram_in_reg_5_4,
	ram_in_reg_6_4,
	ram_in_reg_7_4,
	ram_in_reg_8_4,
	ram_in_reg_4_4,
	ram_in_reg_5_6,
	ram_in_reg_6_6,
	ram_in_reg_7_6,
	ram_in_reg_8_6,
	ram_in_reg_4_6,
	ram_in_reg_3_6,
	ram_in_reg_3_4,
	ram_in_reg_2_6,
	ram_in_reg_2_4,
	ram_in_reg_1_6,
	ram_in_reg_1_4,
	ram_in_reg_0_6,
	ram_in_reg_0_4,
	ram_in_reg_5_5,
	ram_in_reg_6_5,
	ram_in_reg_7_5,
	ram_in_reg_8_5,
	ram_in_reg_4_5,
	ram_in_reg_5_7,
	ram_in_reg_6_7,
	ram_in_reg_7_7,
	ram_in_reg_8_7,
	ram_in_reg_4_7,
	ram_in_reg_3_7,
	ram_in_reg_3_5,
	ram_in_reg_2_7,
	ram_in_reg_2_5,
	ram_in_reg_1_7,
	ram_in_reg_1_5,
	ram_in_reg_0_7,
	ram_in_reg_0_5,
	ram_in_reg_9_4,
	ram_in_reg_9_6,
	ram_in_reg_9_5,
	ram_in_reg_9_7,
	global_clock_enable,
	tdl_arr_0,
	sdetdIDLE,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	Mux1,
	tdl_arr_6,
	reg_no_twiddle605,
	reg_no_twiddle609,
	reg_no_twiddle615,
	reg_no_twiddle619,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_5_12,
	tdl_arr_9_12,
	tdl_arr_5_13,
	tdl_arr_9_13,
	tdl_arr_5_14,
	tdl_arr_9_14,
	tdl_arr_5_15,
	tdl_arr_9_15,
	reg_no_twiddle606,
	reg_no_twiddle616,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	reg_no_twiddle607,
	reg_no_twiddle617,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_7_12,
	tdl_arr_7_13,
	tdl_arr_7_14,
	tdl_arr_7_15,
	reg_no_twiddle608,
	reg_no_twiddle618,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_8_12,
	tdl_arr_8_13,
	tdl_arr_8_14,
	tdl_arr_8_15,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_2_12,
	reg_no_twiddle602,
	tdl_arr_2_13,
	tdl_arr_2_14,
	tdl_arr_2_15,
	reg_no_twiddle612,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_1_12,
	reg_no_twiddle601,
	tdl_arr_1_13,
	tdl_arr_1_14,
	tdl_arr_1_15,
	reg_no_twiddle611,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_0_12,
	reg_no_twiddle600,
	tdl_arr_0_13,
	tdl_arr_0_14,
	tdl_arr_0_15,
	reg_no_twiddle610,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_4_12,
	reg_no_twiddle604,
	tdl_arr_4_13,
	tdl_arr_4_14,
	tdl_arr_4_15,
	reg_no_twiddle614,
	tdl_arr_3_1,
	tdl_arr_3_11,
	tdl_arr_3_12,
	reg_no_twiddle603,
	tdl_arr_3_13,
	tdl_arr_3_14,
	tdl_arr_3_15,
	reg_no_twiddle613,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	ram_in_reg_7_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_8_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_8_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_2_0;
input 	ram_in_reg_1_2;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_8_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_8_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_1;
input 	ram_in_reg_2_3;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_9_0;
input 	ram_in_reg_9_2;
input 	ram_in_reg_9_1;
input 	ram_in_reg_9_3;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_4;
input 	ram_in_reg_8_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_6;
input 	ram_in_reg_8_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_3_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_2_4;
input 	ram_in_reg_1_6;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_5;
input 	ram_in_reg_8_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_8_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_5;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_9_4;
input 	ram_in_reg_9_6;
input 	ram_in_reg_9_5;
input 	ram_in_reg_9_7;
input 	global_clock_enable;
input 	tdl_arr_0;
output 	sdetdIDLE;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	slb_i_0;
output 	slb_i_1;
output 	slb_i_2;
output 	slb_i_3;
output 	Mux2;
output 	Mux1;
input 	tdl_arr_6;
output 	reg_no_twiddle605;
output 	reg_no_twiddle609;
output 	reg_no_twiddle615;
output 	reg_no_twiddle619;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_5_11;
output 	tdl_arr_9_11;
output 	tdl_arr_5_12;
output 	tdl_arr_9_12;
output 	tdl_arr_5_13;
output 	tdl_arr_9_13;
output 	tdl_arr_5_14;
output 	tdl_arr_9_14;
output 	tdl_arr_5_15;
output 	tdl_arr_9_15;
output 	reg_no_twiddle606;
output 	reg_no_twiddle616;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_6_12;
output 	tdl_arr_6_13;
output 	tdl_arr_6_14;
output 	tdl_arr_6_15;
output 	reg_no_twiddle607;
output 	reg_no_twiddle617;
output 	tdl_arr_7_1;
output 	tdl_arr_7_11;
output 	tdl_arr_7_12;
output 	tdl_arr_7_13;
output 	tdl_arr_7_14;
output 	tdl_arr_7_15;
output 	reg_no_twiddle608;
output 	reg_no_twiddle618;
output 	tdl_arr_8_1;
output 	tdl_arr_8_11;
output 	tdl_arr_8_12;
output 	tdl_arr_8_13;
output 	tdl_arr_8_14;
output 	tdl_arr_8_15;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_2_12;
output 	reg_no_twiddle602;
output 	tdl_arr_2_13;
output 	tdl_arr_2_14;
output 	tdl_arr_2_15;
output 	reg_no_twiddle612;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_1_12;
output 	reg_no_twiddle601;
output 	tdl_arr_1_13;
output 	tdl_arr_1_14;
output 	tdl_arr_1_15;
output 	reg_no_twiddle611;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
output 	tdl_arr_0_12;
output 	reg_no_twiddle600;
output 	tdl_arr_0_13;
output 	tdl_arr_0_14;
output 	tdl_arr_0_15;
output 	reg_no_twiddle610;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_4_12;
output 	reg_no_twiddle604;
output 	tdl_arr_4_13;
output 	tdl_arr_4_14;
output 	tdl_arr_4_15;
output 	reg_no_twiddle614;
output 	tdl_arr_3_1;
output 	tdl_arr_3_11;
output 	tdl_arr_3_12;
output 	reg_no_twiddle603;
output 	tdl_arr_3_13;
output 	tdl_arr_3_14;
output 	tdl_arr_3_15;
output 	reg_no_twiddle613;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \butterfly_st2[0][0][8]~q ;
wire \butterfly_st2[0][0][7]~q ;
wire \butterfly_st2[0][0][6]~q ;
wire \butterfly_st2[0][0][5]~q ;
wire \butterfly_st2[0][0][4]~q ;
wire \butterfly_st2[0][0][3]~q ;
wire \butterfly_st2[0][0][2]~q ;
wire \butterfly_st2[0][0][1]~q ;
wire \butterfly_st2[0][0][0]~q ;
wire \butterfly_st2[0][0][11]~q ;
wire \butterfly_st2[0][0][10]~q ;
wire \butterfly_st2[0][0][9]~q ;
wire \butterfly_st2[0][1][8]~q ;
wire \butterfly_st2[0][1][7]~q ;
wire \butterfly_st2[0][1][6]~q ;
wire \butterfly_st2[0][1][5]~q ;
wire \butterfly_st2[0][1][4]~q ;
wire \butterfly_st2[0][1][3]~q ;
wire \butterfly_st2[0][1][2]~q ;
wire \butterfly_st2[0][1][1]~q ;
wire \butterfly_st2[0][1][0]~q ;
wire \butterfly_st2[0][1][11]~q ;
wire \butterfly_st2[0][1][10]~q ;
wire \butterfly_st2[0][1][9]~q ;
wire \butterfly_st2[1][1][2]~q ;
wire \butterfly_st2[1][1][1]~q ;
wire \butterfly_st2[1][1][0]~q ;
wire \butterfly_st2[1][1][11]~q ;
wire \butterfly_st2[1][1][3]~q ;
wire \butterfly_st2[1][1][4]~q ;
wire \butterfly_st2[1][1][5]~q ;
wire \butterfly_st2[1][1][6]~q ;
wire \butterfly_st2[1][1][7]~q ;
wire \butterfly_st2[1][1][8]~q ;
wire \butterfly_st2[1][1][9]~q ;
wire \butterfly_st2[1][1][10]~q ;
wire \butterfly_st2[1][0][2]~q ;
wire \butterfly_st2[1][0][1]~q ;
wire \butterfly_st2[1][0][0]~q ;
wire \butterfly_st2[1][0][11]~q ;
wire \butterfly_st2[1][0][3]~q ;
wire \butterfly_st2[1][0][4]~q ;
wire \butterfly_st2[1][0][5]~q ;
wire \butterfly_st2[1][0][6]~q ;
wire \butterfly_st2[1][0][7]~q ;
wire \butterfly_st2[1][0][8]~q ;
wire \butterfly_st2[1][0][9]~q ;
wire \butterfly_st2[1][0][10]~q ;
wire \butterfly_st2[2][1][2]~q ;
wire \butterfly_st2[2][1][1]~q ;
wire \butterfly_st2[2][1][0]~q ;
wire \butterfly_st2[2][1][11]~q ;
wire \butterfly_st2[2][1][3]~q ;
wire \butterfly_st2[2][1][4]~q ;
wire \butterfly_st2[2][1][5]~q ;
wire \butterfly_st2[2][1][6]~q ;
wire \butterfly_st2[2][1][7]~q ;
wire \butterfly_st2[2][1][8]~q ;
wire \butterfly_st2[2][1][9]~q ;
wire \butterfly_st2[2][1][10]~q ;
wire \butterfly_st2[2][0][2]~q ;
wire \butterfly_st2[2][0][1]~q ;
wire \butterfly_st2[2][0][0]~q ;
wire \butterfly_st2[2][0][11]~q ;
wire \butterfly_st2[2][0][3]~q ;
wire \butterfly_st2[2][0][4]~q ;
wire \butterfly_st2[2][0][5]~q ;
wire \butterfly_st2[2][0][6]~q ;
wire \butterfly_st2[2][0][7]~q ;
wire \butterfly_st2[2][0][8]~q ;
wire \butterfly_st2[2][0][9]~q ;
wire \butterfly_st2[2][0][10]~q ;
wire \butterfly_st2[3][1][2]~q ;
wire \butterfly_st2[3][1][1]~q ;
wire \butterfly_st2[3][1][0]~q ;
wire \butterfly_st2[3][1][11]~q ;
wire \butterfly_st2[3][1][3]~q ;
wire \butterfly_st2[3][1][4]~q ;
wire \butterfly_st2[3][1][5]~q ;
wire \butterfly_st2[3][1][6]~q ;
wire \butterfly_st2[3][1][7]~q ;
wire \butterfly_st2[3][1][8]~q ;
wire \butterfly_st2[3][1][9]~q ;
wire \butterfly_st2[3][1][10]~q ;
wire \butterfly_st2[3][0][2]~q ;
wire \butterfly_st2[3][0][1]~q ;
wire \butterfly_st2[3][0][0]~q ;
wire \butterfly_st2[3][0][11]~q ;
wire \butterfly_st2[3][0][3]~q ;
wire \butterfly_st2[3][0][4]~q ;
wire \butterfly_st2[3][0][5]~q ;
wire \butterfly_st2[3][0][6]~q ;
wire \butterfly_st2[3][0][7]~q ;
wire \butterfly_st2[3][0][8]~q ;
wire \butterfly_st2[3][0][9]~q ;
wire \butterfly_st2[3][0][10]~q ;
wire \butterfly_st1[0][0][8]~q ;
wire \butterfly_st1[1][0][8]~q ;
wire \butterfly_st1[0][0][7]~q ;
wire \butterfly_st1[1][0][7]~q ;
wire \butterfly_st1[0][0][6]~q ;
wire \butterfly_st1[1][0][6]~q ;
wire \butterfly_st1[0][0][5]~q ;
wire \butterfly_st1[1][0][5]~q ;
wire \butterfly_st1[0][0][4]~q ;
wire \butterfly_st1[1][0][4]~q ;
wire \butterfly_st1[0][0][3]~q ;
wire \butterfly_st1[1][0][3]~q ;
wire \butterfly_st1[0][0][2]~q ;
wire \butterfly_st1[1][0][2]~q ;
wire \butterfly_st1[0][0][1]~q ;
wire \butterfly_st1[1][0][1]~q ;
wire \butterfly_st1[0][0][0]~q ;
wire \butterfly_st1[1][0][0]~q ;
wire \butterfly_st2[0][0][0]~2 ;
wire \butterfly_st2[0][0][0]~1_combout ;
wire \butterfly_st2[0][0][1]~2 ;
wire \butterfly_st2[0][0][1]~1_combout ;
wire \butterfly_st2[0][0][2]~2 ;
wire \butterfly_st2[0][0][2]~1_combout ;
wire \butterfly_st2[0][0][3]~2 ;
wire \butterfly_st2[0][0][3]~1_combout ;
wire \butterfly_st2[0][0][4]~2 ;
wire \butterfly_st2[0][0][4]~1_combout ;
wire \butterfly_st2[0][0][5]~2 ;
wire \butterfly_st2[0][0][5]~1_combout ;
wire \butterfly_st2[0][0][6]~2 ;
wire \butterfly_st2[0][0][6]~1_combout ;
wire \butterfly_st2[0][0][7]~2 ;
wire \butterfly_st2[0][0][7]~1_combout ;
wire \butterfly_st2[0][0][8]~2 ;
wire \butterfly_st2[0][0][8]~1_combout ;
wire \butterfly_st1[0][0][10]~q ;
wire \butterfly_st1[1][0][10]~q ;
wire \butterfly_st1[0][0][9]~q ;
wire \butterfly_st1[1][0][9]~q ;
wire \butterfly_st2[0][0][9]~2 ;
wire \butterfly_st2[0][0][9]~1_combout ;
wire \butterfly_st2[0][0][10]~2 ;
wire \butterfly_st2[0][0][10]~1_combout ;
wire \butterfly_st2[0][0][11]~1_combout ;
wire \butterfly_st1[0][1][8]~q ;
wire \butterfly_st1[1][1][8]~q ;
wire \butterfly_st1[0][1][7]~q ;
wire \butterfly_st1[1][1][7]~q ;
wire \butterfly_st1[0][1][6]~q ;
wire \butterfly_st1[1][1][6]~q ;
wire \butterfly_st1[0][1][5]~q ;
wire \butterfly_st1[1][1][5]~q ;
wire \butterfly_st1[0][1][4]~q ;
wire \butterfly_st1[1][1][4]~q ;
wire \butterfly_st1[0][1][3]~q ;
wire \butterfly_st1[1][1][3]~q ;
wire \butterfly_st1[0][1][2]~q ;
wire \butterfly_st1[1][1][2]~q ;
wire \butterfly_st1[0][1][1]~q ;
wire \butterfly_st1[1][1][1]~q ;
wire \butterfly_st1[0][1][0]~q ;
wire \butterfly_st1[1][1][0]~q ;
wire \butterfly_st2[0][1][0]~2 ;
wire \butterfly_st2[0][1][0]~1_combout ;
wire \butterfly_st2[0][1][1]~2 ;
wire \butterfly_st2[0][1][1]~1_combout ;
wire \butterfly_st2[0][1][2]~2 ;
wire \butterfly_st2[0][1][2]~1_combout ;
wire \butterfly_st2[0][1][3]~2 ;
wire \butterfly_st2[0][1][3]~1_combout ;
wire \butterfly_st2[0][1][4]~2 ;
wire \butterfly_st2[0][1][4]~1_combout ;
wire \butterfly_st2[0][1][5]~2 ;
wire \butterfly_st2[0][1][5]~1_combout ;
wire \butterfly_st2[0][1][6]~2 ;
wire \butterfly_st2[0][1][6]~1_combout ;
wire \butterfly_st2[0][1][7]~2 ;
wire \butterfly_st2[0][1][7]~1_combout ;
wire \butterfly_st2[0][1][8]~2 ;
wire \butterfly_st2[0][1][8]~1_combout ;
wire \butterfly_st1[0][1][10]~q ;
wire \butterfly_st1[1][1][10]~q ;
wire \butterfly_st1[0][1][9]~q ;
wire \butterfly_st1[1][1][9]~q ;
wire \butterfly_st2[0][1][9]~2 ;
wire \butterfly_st2[0][1][9]~1_combout ;
wire \butterfly_st2[0][1][10]~2 ;
wire \butterfly_st2[0][1][10]~1_combout ;
wire \butterfly_st2[0][1][11]~1_combout ;
wire \butterfly_st1[2][1][2]~q ;
wire \butterfly_st1[3][0][2]~q ;
wire \butterfly_st1[2][1][1]~q ;
wire \butterfly_st1[3][0][1]~q ;
wire \butterfly_st1[2][1][0]~q ;
wire \butterfly_st1[3][0][0]~q ;
wire \butterfly_st2[1][1][0]~2 ;
wire \butterfly_st2[1][1][0]~1_combout ;
wire \butterfly_st2[1][1][1]~2 ;
wire \butterfly_st2[1][1][1]~1_combout ;
wire \butterfly_st2[1][1][2]~2 ;
wire \butterfly_st2[1][1][2]~1_combout ;
wire \butterfly_st1[2][1][10]~q ;
wire \butterfly_st1[3][0][10]~q ;
wire \butterfly_st1[2][1][9]~q ;
wire \butterfly_st1[3][0][9]~q ;
wire \butterfly_st1[2][1][8]~q ;
wire \butterfly_st1[3][0][8]~q ;
wire \butterfly_st1[2][1][7]~q ;
wire \butterfly_st1[3][0][7]~q ;
wire \butterfly_st1[2][1][6]~q ;
wire \butterfly_st1[3][0][6]~q ;
wire \butterfly_st1[2][1][5]~q ;
wire \butterfly_st1[3][0][5]~q ;
wire \butterfly_st1[2][1][4]~q ;
wire \butterfly_st1[3][0][4]~q ;
wire \butterfly_st1[2][1][3]~q ;
wire \butterfly_st1[3][0][3]~q ;
wire \butterfly_st2[1][1][3]~2 ;
wire \butterfly_st2[1][1][3]~1_combout ;
wire \butterfly_st2[1][1][4]~2 ;
wire \butterfly_st2[1][1][4]~1_combout ;
wire \butterfly_st2[1][1][5]~2 ;
wire \butterfly_st2[1][1][5]~1_combout ;
wire \butterfly_st2[1][1][6]~2 ;
wire \butterfly_st2[1][1][6]~1_combout ;
wire \butterfly_st2[1][1][7]~2 ;
wire \butterfly_st2[1][1][7]~1_combout ;
wire \butterfly_st2[1][1][8]~2 ;
wire \butterfly_st2[1][1][8]~1_combout ;
wire \butterfly_st2[1][1][9]~2 ;
wire \butterfly_st2[1][1][9]~1_combout ;
wire \butterfly_st2[1][1][10]~2 ;
wire \butterfly_st2[1][1][10]~1_combout ;
wire \butterfly_st2[1][1][11]~1_combout ;
wire \butterfly_st1[2][0][2]~q ;
wire \butterfly_st1[3][1][2]~q ;
wire \butterfly_st1[2][0][1]~q ;
wire \butterfly_st1[3][1][1]~q ;
wire \butterfly_st1[2][0][0]~q ;
wire \butterfly_st1[3][1][0]~q ;
wire \butterfly_st2[1][0][0]~2 ;
wire \butterfly_st2[1][0][0]~1_combout ;
wire \butterfly_st2[1][0][1]~2 ;
wire \butterfly_st2[1][0][1]~1_combout ;
wire \butterfly_st2[1][0][2]~2 ;
wire \butterfly_st2[1][0][2]~1_combout ;
wire \butterfly_st1[2][0][10]~q ;
wire \butterfly_st1[3][1][10]~q ;
wire \butterfly_st1[2][0][9]~q ;
wire \butterfly_st1[3][1][9]~q ;
wire \butterfly_st1[2][0][8]~q ;
wire \butterfly_st1[3][1][8]~q ;
wire \butterfly_st1[2][0][7]~q ;
wire \butterfly_st1[3][1][7]~q ;
wire \butterfly_st1[2][0][6]~q ;
wire \butterfly_st1[3][1][6]~q ;
wire \butterfly_st1[2][0][5]~q ;
wire \butterfly_st1[3][1][5]~q ;
wire \butterfly_st1[2][0][4]~q ;
wire \butterfly_st1[3][1][4]~q ;
wire \butterfly_st1[2][0][3]~q ;
wire \butterfly_st1[3][1][3]~q ;
wire \butterfly_st2[1][0][3]~2 ;
wire \butterfly_st2[1][0][3]~1_combout ;
wire \butterfly_st2[1][0][4]~2 ;
wire \butterfly_st2[1][0][4]~1_combout ;
wire \butterfly_st2[1][0][5]~2 ;
wire \butterfly_st2[1][0][5]~1_combout ;
wire \butterfly_st2[1][0][6]~2 ;
wire \butterfly_st2[1][0][6]~1_combout ;
wire \butterfly_st2[1][0][7]~2 ;
wire \butterfly_st2[1][0][7]~1_combout ;
wire \butterfly_st2[1][0][8]~2 ;
wire \butterfly_st2[1][0][8]~1_combout ;
wire \butterfly_st2[1][0][9]~2 ;
wire \butterfly_st2[1][0][9]~1_combout ;
wire \butterfly_st2[1][0][10]~2 ;
wire \butterfly_st2[1][0][10]~1_combout ;
wire \butterfly_st2[1][0][11]~1_combout ;
wire \butterfly_st2[2][1][0]~2 ;
wire \butterfly_st2[2][1][0]~1_combout ;
wire \butterfly_st2[2][1][1]~2 ;
wire \butterfly_st2[2][1][1]~1_combout ;
wire \butterfly_st2[2][1][2]~2 ;
wire \butterfly_st2[2][1][2]~1_combout ;
wire \butterfly_st2[2][1][3]~2 ;
wire \butterfly_st2[2][1][3]~1_combout ;
wire \butterfly_st2[2][1][4]~2 ;
wire \butterfly_st2[2][1][4]~1_combout ;
wire \butterfly_st2[2][1][5]~2 ;
wire \butterfly_st2[2][1][5]~1_combout ;
wire \butterfly_st2[2][1][6]~2 ;
wire \butterfly_st2[2][1][6]~1_combout ;
wire \butterfly_st2[2][1][7]~2 ;
wire \butterfly_st2[2][1][7]~1_combout ;
wire \butterfly_st2[2][1][8]~2 ;
wire \butterfly_st2[2][1][8]~1_combout ;
wire \butterfly_st2[2][1][9]~2 ;
wire \butterfly_st2[2][1][9]~1_combout ;
wire \butterfly_st2[2][1][10]~2 ;
wire \butterfly_st2[2][1][10]~1_combout ;
wire \butterfly_st2[2][1][11]~1_combout ;
wire \butterfly_st2[2][0][0]~2 ;
wire \butterfly_st2[2][0][0]~1_combout ;
wire \butterfly_st2[2][0][1]~2 ;
wire \butterfly_st2[2][0][1]~1_combout ;
wire \butterfly_st2[2][0][2]~2 ;
wire \butterfly_st2[2][0][2]~1_combout ;
wire \butterfly_st2[2][0][3]~2 ;
wire \butterfly_st2[2][0][3]~1_combout ;
wire \butterfly_st2[2][0][4]~2 ;
wire \butterfly_st2[2][0][4]~1_combout ;
wire \butterfly_st2[2][0][5]~2 ;
wire \butterfly_st2[2][0][5]~1_combout ;
wire \butterfly_st2[2][0][6]~2 ;
wire \butterfly_st2[2][0][6]~1_combout ;
wire \butterfly_st2[2][0][7]~2 ;
wire \butterfly_st2[2][0][7]~1_combout ;
wire \butterfly_st2[2][0][8]~2 ;
wire \butterfly_st2[2][0][8]~1_combout ;
wire \butterfly_st2[2][0][9]~2 ;
wire \butterfly_st2[2][0][9]~1_combout ;
wire \butterfly_st2[2][0][10]~2 ;
wire \butterfly_st2[2][0][10]~1_combout ;
wire \butterfly_st2[2][0][11]~1_combout ;
wire \butterfly_st2[3][1][0]~2 ;
wire \butterfly_st2[3][1][0]~1_combout ;
wire \butterfly_st2[3][1][1]~2 ;
wire \butterfly_st2[3][1][1]~1_combout ;
wire \butterfly_st2[3][1][2]~2 ;
wire \butterfly_st2[3][1][2]~1_combout ;
wire \butterfly_st2[3][1][3]~2 ;
wire \butterfly_st2[3][1][3]~1_combout ;
wire \butterfly_st2[3][1][4]~2 ;
wire \butterfly_st2[3][1][4]~1_combout ;
wire \butterfly_st2[3][1][5]~2 ;
wire \butterfly_st2[3][1][5]~1_combout ;
wire \butterfly_st2[3][1][6]~2 ;
wire \butterfly_st2[3][1][6]~1_combout ;
wire \butterfly_st2[3][1][7]~2 ;
wire \butterfly_st2[3][1][7]~1_combout ;
wire \butterfly_st2[3][1][8]~2 ;
wire \butterfly_st2[3][1][8]~1_combout ;
wire \butterfly_st2[3][1][9]~2 ;
wire \butterfly_st2[3][1][9]~1_combout ;
wire \butterfly_st2[3][1][10]~2 ;
wire \butterfly_st2[3][1][10]~1_combout ;
wire \butterfly_st2[3][1][11]~1_combout ;
wire \butterfly_st2[3][0][0]~2 ;
wire \butterfly_st2[3][0][0]~1_combout ;
wire \butterfly_st2[3][0][1]~2 ;
wire \butterfly_st2[3][0][1]~1_combout ;
wire \butterfly_st2[3][0][2]~2 ;
wire \butterfly_st2[3][0][2]~1_combout ;
wire \butterfly_st2[3][0][3]~2 ;
wire \butterfly_st2[3][0][3]~1_combout ;
wire \butterfly_st2[3][0][4]~2 ;
wire \butterfly_st2[3][0][4]~1_combout ;
wire \butterfly_st2[3][0][5]~2 ;
wire \butterfly_st2[3][0][5]~1_combout ;
wire \butterfly_st2[3][0][6]~2 ;
wire \butterfly_st2[3][0][6]~1_combout ;
wire \butterfly_st2[3][0][7]~2 ;
wire \butterfly_st2[3][0][7]~1_combout ;
wire \butterfly_st2[3][0][8]~2 ;
wire \butterfly_st2[3][0][8]~1_combout ;
wire \butterfly_st2[3][0][9]~2 ;
wire \butterfly_st2[3][0][9]~1_combout ;
wire \butterfly_st2[3][0][10]~2 ;
wire \butterfly_st2[3][0][10]~1_combout ;
wire \butterfly_st2[3][0][11]~1_combout ;
wire \gen_disc:bfp_scale|r_array_out[2][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][2]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][2]~q ;
wire \butterfly_st1[0][0][0]~2 ;
wire \butterfly_st1[0][0][0]~1_combout ;
wire \butterfly_st1[0][0][1]~2 ;
wire \butterfly_st1[0][0][1]~1_combout ;
wire \butterfly_st1[0][0][2]~2 ;
wire \butterfly_st1[0][0][2]~1_combout ;
wire \butterfly_st1[0][0][3]~2 ;
wire \butterfly_st1[0][0][3]~1_combout ;
wire \butterfly_st1[0][0][4]~2 ;
wire \butterfly_st1[0][0][4]~1_combout ;
wire \butterfly_st1[0][0][5]~2 ;
wire \butterfly_st1[0][0][5]~1_combout ;
wire \butterfly_st1[0][0][6]~2 ;
wire \butterfly_st1[0][0][6]~1_combout ;
wire \butterfly_st1[0][0][7]~2 ;
wire \butterfly_st1[0][0][7]~1_combout ;
wire \butterfly_st1[0][0][8]~2 ;
wire \butterfly_st1[0][0][8]~1_combout ;
wire \gen_disc:bfp_scale|r_array_out[3][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][2]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][2]~q ;
wire \butterfly_st1[1][0][0]~2 ;
wire \butterfly_st1[1][0][0]~1_combout ;
wire \butterfly_st1[1][0][1]~2 ;
wire \butterfly_st1[1][0][1]~1_combout ;
wire \butterfly_st1[1][0][2]~2 ;
wire \butterfly_st1[1][0][2]~1_combout ;
wire \butterfly_st1[1][0][3]~2 ;
wire \butterfly_st1[1][0][3]~1_combout ;
wire \butterfly_st1[1][0][4]~2 ;
wire \butterfly_st1[1][0][4]~1_combout ;
wire \butterfly_st1[1][0][5]~2 ;
wire \butterfly_st1[1][0][5]~1_combout ;
wire \butterfly_st1[1][0][6]~2 ;
wire \butterfly_st1[1][0][6]~1_combout ;
wire \butterfly_st1[1][0][7]~2 ;
wire \butterfly_st1[1][0][7]~1_combout ;
wire \butterfly_st1[1][0][8]~2 ;
wire \butterfly_st1[1][0][8]~1_combout ;
wire \butterfly_st1[0][0][9]~2 ;
wire \butterfly_st1[0][0][9]~1_combout ;
wire \butterfly_st1[0][0][10]~1_combout ;
wire \butterfly_st1[1][0][9]~2 ;
wire \butterfly_st1[1][0][9]~1_combout ;
wire \butterfly_st1[1][0][10]~1_combout ;
wire \gen_disc:bfp_scale|i_array_out[2][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][2]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][2]~q ;
wire \butterfly_st1[0][1][0]~2 ;
wire \butterfly_st1[0][1][0]~1_combout ;
wire \butterfly_st1[0][1][1]~2 ;
wire \butterfly_st1[0][1][1]~1_combout ;
wire \butterfly_st1[0][1][2]~2 ;
wire \butterfly_st1[0][1][2]~1_combout ;
wire \butterfly_st1[0][1][3]~2 ;
wire \butterfly_st1[0][1][3]~1_combout ;
wire \butterfly_st1[0][1][4]~2 ;
wire \butterfly_st1[0][1][4]~1_combout ;
wire \butterfly_st1[0][1][5]~2 ;
wire \butterfly_st1[0][1][5]~1_combout ;
wire \butterfly_st1[0][1][6]~2 ;
wire \butterfly_st1[0][1][6]~1_combout ;
wire \butterfly_st1[0][1][7]~2 ;
wire \butterfly_st1[0][1][7]~1_combout ;
wire \butterfly_st1[0][1][8]~2 ;
wire \butterfly_st1[0][1][8]~1_combout ;
wire \gen_disc:bfp_scale|i_array_out[3][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][2]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][2]~q ;
wire \butterfly_st1[1][1][0]~2 ;
wire \butterfly_st1[1][1][0]~1_combout ;
wire \butterfly_st1[1][1][1]~2 ;
wire \butterfly_st1[1][1][1]~1_combout ;
wire \butterfly_st1[1][1][2]~2 ;
wire \butterfly_st1[1][1][2]~1_combout ;
wire \butterfly_st1[1][1][3]~2 ;
wire \butterfly_st1[1][1][3]~1_combout ;
wire \butterfly_st1[1][1][4]~2 ;
wire \butterfly_st1[1][1][4]~1_combout ;
wire \butterfly_st1[1][1][5]~2 ;
wire \butterfly_st1[1][1][5]~1_combout ;
wire \butterfly_st1[1][1][6]~2 ;
wire \butterfly_st1[1][1][6]~1_combout ;
wire \butterfly_st1[1][1][7]~2 ;
wire \butterfly_st1[1][1][7]~1_combout ;
wire \butterfly_st1[1][1][8]~2 ;
wire \butterfly_st1[1][1][8]~1_combout ;
wire \butterfly_st1[0][1][9]~2 ;
wire \butterfly_st1[0][1][9]~1_combout ;
wire \butterfly_st1[0][1][10]~1_combout ;
wire \butterfly_st1[1][1][9]~2 ;
wire \butterfly_st1[1][1][9]~1_combout ;
wire \butterfly_st1[1][1][10]~1_combout ;
wire \butterfly_st1[2][1][0]~2 ;
wire \butterfly_st1[2][1][0]~1_combout ;
wire \butterfly_st1[2][1][1]~2 ;
wire \butterfly_st1[2][1][1]~1_combout ;
wire \butterfly_st1[2][1][2]~2 ;
wire \butterfly_st1[2][1][2]~1_combout ;
wire \butterfly_st1[3][0][0]~2 ;
wire \butterfly_st1[3][0][0]~1_combout ;
wire \butterfly_st1[3][0][1]~2 ;
wire \butterfly_st1[3][0][1]~1_combout ;
wire \butterfly_st1[3][0][2]~2 ;
wire \butterfly_st1[3][0][2]~1_combout ;
wire \butterfly_st1[2][1][3]~2 ;
wire \butterfly_st1[2][1][3]~1_combout ;
wire \butterfly_st1[2][1][4]~2 ;
wire \butterfly_st1[2][1][4]~1_combout ;
wire \butterfly_st1[2][1][5]~2 ;
wire \butterfly_st1[2][1][5]~1_combout ;
wire \butterfly_st1[2][1][6]~2 ;
wire \butterfly_st1[2][1][6]~1_combout ;
wire \butterfly_st1[2][1][7]~2 ;
wire \butterfly_st1[2][1][7]~1_combout ;
wire \butterfly_st1[2][1][8]~2 ;
wire \butterfly_st1[2][1][8]~1_combout ;
wire \butterfly_st1[2][1][9]~2 ;
wire \butterfly_st1[2][1][9]~1_combout ;
wire \butterfly_st1[2][1][10]~1_combout ;
wire \butterfly_st1[3][0][3]~2 ;
wire \butterfly_st1[3][0][3]~1_combout ;
wire \butterfly_st1[3][0][4]~2 ;
wire \butterfly_st1[3][0][4]~1_combout ;
wire \butterfly_st1[3][0][5]~2 ;
wire \butterfly_st1[3][0][5]~1_combout ;
wire \butterfly_st1[3][0][6]~2 ;
wire \butterfly_st1[3][0][6]~1_combout ;
wire \butterfly_st1[3][0][7]~2 ;
wire \butterfly_st1[3][0][7]~1_combout ;
wire \butterfly_st1[3][0][8]~2 ;
wire \butterfly_st1[3][0][8]~1_combout ;
wire \butterfly_st1[3][0][9]~2 ;
wire \butterfly_st1[3][0][9]~1_combout ;
wire \butterfly_st1[3][0][10]~1_combout ;
wire \butterfly_st1[2][0][0]~2 ;
wire \butterfly_st1[2][0][0]~1_combout ;
wire \butterfly_st1[2][0][1]~2 ;
wire \butterfly_st1[2][0][1]~1_combout ;
wire \butterfly_st1[2][0][2]~2 ;
wire \butterfly_st1[2][0][2]~1_combout ;
wire \butterfly_st1[3][1][0]~2 ;
wire \butterfly_st1[3][1][0]~1_combout ;
wire \butterfly_st1[3][1][1]~2 ;
wire \butterfly_st1[3][1][1]~1_combout ;
wire \butterfly_st1[3][1][2]~2 ;
wire \butterfly_st1[3][1][2]~1_combout ;
wire \butterfly_st1[2][0][3]~2 ;
wire \butterfly_st1[2][0][3]~1_combout ;
wire \butterfly_st1[2][0][4]~2 ;
wire \butterfly_st1[2][0][4]~1_combout ;
wire \butterfly_st1[2][0][5]~2 ;
wire \butterfly_st1[2][0][5]~1_combout ;
wire \butterfly_st1[2][0][6]~2 ;
wire \butterfly_st1[2][0][6]~1_combout ;
wire \butterfly_st1[2][0][7]~2 ;
wire \butterfly_st1[2][0][7]~1_combout ;
wire \butterfly_st1[2][0][8]~2 ;
wire \butterfly_st1[2][0][8]~1_combout ;
wire \butterfly_st1[2][0][9]~2 ;
wire \butterfly_st1[2][0][9]~1_combout ;
wire \butterfly_st1[2][0][10]~1_combout ;
wire \butterfly_st1[3][1][3]~2 ;
wire \butterfly_st1[3][1][3]~1_combout ;
wire \butterfly_st1[3][1][4]~2 ;
wire \butterfly_st1[3][1][4]~1_combout ;
wire \butterfly_st1[3][1][5]~2 ;
wire \butterfly_st1[3][1][5]~1_combout ;
wire \butterfly_st1[3][1][6]~2 ;
wire \butterfly_st1[3][1][6]~1_combout ;
wire \butterfly_st1[3][1][7]~2 ;
wire \butterfly_st1[3][1][7]~1_combout ;
wire \butterfly_st1[3][1][8]~2 ;
wire \butterfly_st1[3][1][8]~1_combout ;
wire \butterfly_st1[3][1][9]~2 ;
wire \butterfly_st1[3][1][9]~1_combout ;
wire \butterfly_st1[3][1][10]~1_combout ;
wire \gen_disc:bfp_scale|r_array_out[0][8]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][8]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][8]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][8]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][9]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][9]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][9]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][9]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][8]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][8]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][8]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][8]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][9]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][9]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][9]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][9]~q ;
wire \reg_no_twiddle~80_combout ;
wire \reg_no_twiddle[0][0][0]~2 ;
wire \reg_no_twiddle[0][0][1]~2 ;
wire \reg_no_twiddle[0][0][2]~2 ;
wire \reg_no_twiddle[0][0][3]~2 ;
wire \reg_no_twiddle[0][0][4]~2 ;
wire \reg_no_twiddle[0][0][5]~1_combout ;
wire \reg_no_twiddle[0][0][5]~q ;
wire \reg_no_twiddle~60_combout ;
wire \reg_no_twiddle[1][0][5]~q ;
wire \reg_no_twiddle~40_combout ;
wire \reg_no_twiddle[2][0][5]~q ;
wire \reg_no_twiddle~30_combout ;
wire \reg_no_twiddle[3][0][5]~q ;
wire \reg_no_twiddle~20_combout ;
wire \reg_no_twiddle[4][0][5]~q ;
wire \reg_no_twiddle~10_combout ;
wire \reg_no_twiddle[5][0][5]~q ;
wire \reg_no_twiddle~0_combout ;
wire \reg_no_twiddle[0][0][5]~2 ;
wire \reg_no_twiddle[0][0][6]~2 ;
wire \reg_no_twiddle[0][0][7]~2 ;
wire \reg_no_twiddle[0][0][8]~2 ;
wire \reg_no_twiddle[0][0][9]~1_combout ;
wire \reg_no_twiddle[0][0][9]~q ;
wire \reg_no_twiddle~61_combout ;
wire \reg_no_twiddle[1][0][9]~q ;
wire \reg_no_twiddle~41_combout ;
wire \reg_no_twiddle[2][0][9]~q ;
wire \reg_no_twiddle~31_combout ;
wire \reg_no_twiddle[3][0][9]~q ;
wire \reg_no_twiddle~21_combout ;
wire \reg_no_twiddle[4][0][9]~q ;
wire \reg_no_twiddle~11_combout ;
wire \reg_no_twiddle[5][0][9]~q ;
wire \reg_no_twiddle~1_combout ;
wire \reg_no_twiddle~81_combout ;
wire \reg_no_twiddle[0][1][0]~2 ;
wire \reg_no_twiddle[0][1][1]~2 ;
wire \reg_no_twiddle[0][1][2]~2 ;
wire \reg_no_twiddle[0][1][3]~2 ;
wire \reg_no_twiddle[0][1][4]~2 ;
wire \reg_no_twiddle[0][1][5]~1_combout ;
wire \reg_no_twiddle[0][1][5]~q ;
wire \reg_no_twiddle~62_combout ;
wire \reg_no_twiddle[1][1][5]~q ;
wire \reg_no_twiddle~42_combout ;
wire \reg_no_twiddle[2][1][5]~q ;
wire \reg_no_twiddle~32_combout ;
wire \reg_no_twiddle[3][1][5]~q ;
wire \reg_no_twiddle~22_combout ;
wire \reg_no_twiddle[4][1][5]~q ;
wire \reg_no_twiddle~12_combout ;
wire \reg_no_twiddle[5][1][5]~q ;
wire \reg_no_twiddle~2_combout ;
wire \reg_no_twiddle[0][1][5]~2 ;
wire \reg_no_twiddle[0][1][6]~2 ;
wire \reg_no_twiddle[0][1][7]~2 ;
wire \reg_no_twiddle[0][1][8]~2 ;
wire \reg_no_twiddle[0][1][9]~1_combout ;
wire \reg_no_twiddle[0][1][9]~q ;
wire \reg_no_twiddle~63_combout ;
wire \reg_no_twiddle[1][1][9]~q ;
wire \reg_no_twiddle~43_combout ;
wire \reg_no_twiddle[2][1][9]~q ;
wire \reg_no_twiddle~33_combout ;
wire \reg_no_twiddle[3][1][9]~q ;
wire \reg_no_twiddle~23_combout ;
wire \reg_no_twiddle[4][1][9]~q ;
wire \reg_no_twiddle~13_combout ;
wire \reg_no_twiddle[5][1][9]~q ;
wire \reg_no_twiddle~3_combout ;
wire \reg_no_twiddle[0][0][6]~1_combout ;
wire \reg_no_twiddle[0][0][6]~q ;
wire \reg_no_twiddle~64_combout ;
wire \reg_no_twiddle[1][0][6]~q ;
wire \reg_no_twiddle~44_combout ;
wire \reg_no_twiddle[2][0][6]~q ;
wire \reg_no_twiddle~34_combout ;
wire \reg_no_twiddle[3][0][6]~q ;
wire \reg_no_twiddle~24_combout ;
wire \reg_no_twiddle[4][0][6]~q ;
wire \reg_no_twiddle~14_combout ;
wire \reg_no_twiddle[5][0][6]~q ;
wire \reg_no_twiddle~4_combout ;
wire \reg_no_twiddle[0][1][6]~1_combout ;
wire \reg_no_twiddle[0][1][6]~q ;
wire \reg_no_twiddle~65_combout ;
wire \reg_no_twiddle[1][1][6]~q ;
wire \reg_no_twiddle~45_combout ;
wire \reg_no_twiddle[2][1][6]~q ;
wire \reg_no_twiddle~35_combout ;
wire \reg_no_twiddle[3][1][6]~q ;
wire \reg_no_twiddle~25_combout ;
wire \reg_no_twiddle[4][1][6]~q ;
wire \reg_no_twiddle~15_combout ;
wire \reg_no_twiddle[5][1][6]~q ;
wire \reg_no_twiddle~5_combout ;
wire \reg_no_twiddle[0][0][7]~1_combout ;
wire \reg_no_twiddle[0][0][7]~q ;
wire \reg_no_twiddle~66_combout ;
wire \reg_no_twiddle[1][0][7]~q ;
wire \reg_no_twiddle~46_combout ;
wire \reg_no_twiddle[2][0][7]~q ;
wire \reg_no_twiddle~36_combout ;
wire \reg_no_twiddle[3][0][7]~q ;
wire \reg_no_twiddle~26_combout ;
wire \reg_no_twiddle[4][0][7]~q ;
wire \reg_no_twiddle~16_combout ;
wire \reg_no_twiddle[5][0][7]~q ;
wire \reg_no_twiddle~6_combout ;
wire \reg_no_twiddle[0][1][7]~1_combout ;
wire \reg_no_twiddle[0][1][7]~q ;
wire \reg_no_twiddle~67_combout ;
wire \reg_no_twiddle[1][1][7]~q ;
wire \reg_no_twiddle~47_combout ;
wire \reg_no_twiddle[2][1][7]~q ;
wire \reg_no_twiddle~37_combout ;
wire \reg_no_twiddle[3][1][7]~q ;
wire \reg_no_twiddle~27_combout ;
wire \reg_no_twiddle[4][1][7]~q ;
wire \reg_no_twiddle~17_combout ;
wire \reg_no_twiddle[5][1][7]~q ;
wire \reg_no_twiddle~7_combout ;
wire \reg_no_twiddle[0][0][8]~1_combout ;
wire \reg_no_twiddle[0][0][8]~q ;
wire \reg_no_twiddle~68_combout ;
wire \reg_no_twiddle[1][0][8]~q ;
wire \reg_no_twiddle~48_combout ;
wire \reg_no_twiddle[2][0][8]~q ;
wire \reg_no_twiddle~38_combout ;
wire \reg_no_twiddle[3][0][8]~q ;
wire \reg_no_twiddle~28_combout ;
wire \reg_no_twiddle[4][0][8]~q ;
wire \reg_no_twiddle~18_combout ;
wire \reg_no_twiddle[5][0][8]~q ;
wire \reg_no_twiddle~8_combout ;
wire \reg_no_twiddle[0][1][8]~1_combout ;
wire \reg_no_twiddle[0][1][8]~q ;
wire \reg_no_twiddle~69_combout ;
wire \reg_no_twiddle[1][1][8]~q ;
wire \reg_no_twiddle~49_combout ;
wire \reg_no_twiddle[2][1][8]~q ;
wire \reg_no_twiddle~39_combout ;
wire \reg_no_twiddle[3][1][8]~q ;
wire \reg_no_twiddle~29_combout ;
wire \reg_no_twiddle[4][1][8]~q ;
wire \reg_no_twiddle~19_combout ;
wire \reg_no_twiddle[5][1][8]~q ;
wire \reg_no_twiddle~9_combout ;
wire \reg_no_twiddle[0][0][2]~1_combout ;
wire \reg_no_twiddle[0][0][2]~q ;
wire \reg_no_twiddle~112_combout ;
wire \reg_no_twiddle[1][0][2]~q ;
wire \reg_no_twiddle~102_combout ;
wire \reg_no_twiddle[2][0][2]~q ;
wire \reg_no_twiddle~92_combout ;
wire \reg_no_twiddle[3][0][2]~q ;
wire \reg_no_twiddle~82_combout ;
wire \reg_no_twiddle[4][0][2]~q ;
wire \reg_no_twiddle~70_combout ;
wire \reg_no_twiddle[5][0][2]~q ;
wire \reg_no_twiddle~50_combout ;
wire \reg_no_twiddle[0][1][2]~1_combout ;
wire \reg_no_twiddle[0][1][2]~q ;
wire \reg_no_twiddle~113_combout ;
wire \reg_no_twiddle[1][1][2]~q ;
wire \reg_no_twiddle~103_combout ;
wire \reg_no_twiddle[2][1][2]~q ;
wire \reg_no_twiddle~93_combout ;
wire \reg_no_twiddle[3][1][2]~q ;
wire \reg_no_twiddle~83_combout ;
wire \reg_no_twiddle[4][1][2]~q ;
wire \reg_no_twiddle~71_combout ;
wire \reg_no_twiddle[5][1][2]~q ;
wire \reg_no_twiddle~51_combout ;
wire \reg_no_twiddle[0][0][1]~1_combout ;
wire \reg_no_twiddle[0][0][1]~q ;
wire \reg_no_twiddle~114_combout ;
wire \reg_no_twiddle[1][0][1]~q ;
wire \reg_no_twiddle~104_combout ;
wire \reg_no_twiddle[2][0][1]~q ;
wire \reg_no_twiddle~94_combout ;
wire \reg_no_twiddle[3][0][1]~q ;
wire \reg_no_twiddle~84_combout ;
wire \reg_no_twiddle[4][0][1]~q ;
wire \reg_no_twiddle~72_combout ;
wire \reg_no_twiddle[5][0][1]~q ;
wire \reg_no_twiddle~52_combout ;
wire \reg_no_twiddle[0][1][1]~1_combout ;
wire \reg_no_twiddle[0][1][1]~q ;
wire \reg_no_twiddle~115_combout ;
wire \reg_no_twiddle[1][1][1]~q ;
wire \reg_no_twiddle~105_combout ;
wire \reg_no_twiddle[2][1][1]~q ;
wire \reg_no_twiddle~95_combout ;
wire \reg_no_twiddle[3][1][1]~q ;
wire \reg_no_twiddle~85_combout ;
wire \reg_no_twiddle[4][1][1]~q ;
wire \reg_no_twiddle~73_combout ;
wire \reg_no_twiddle[5][1][1]~q ;
wire \reg_no_twiddle~53_combout ;
wire \reg_no_twiddle[0][0][0]~1_combout ;
wire \reg_no_twiddle[0][0][0]~q ;
wire \reg_no_twiddle~116_combout ;
wire \reg_no_twiddle[1][0][0]~q ;
wire \reg_no_twiddle~106_combout ;
wire \reg_no_twiddle[2][0][0]~q ;
wire \reg_no_twiddle~96_combout ;
wire \reg_no_twiddle[3][0][0]~q ;
wire \reg_no_twiddle~86_combout ;
wire \reg_no_twiddle[4][0][0]~q ;
wire \reg_no_twiddle~74_combout ;
wire \reg_no_twiddle[5][0][0]~q ;
wire \reg_no_twiddle~54_combout ;
wire \reg_no_twiddle[0][1][0]~1_combout ;
wire \reg_no_twiddle[0][1][0]~q ;
wire \reg_no_twiddle~117_combout ;
wire \reg_no_twiddle[1][1][0]~q ;
wire \reg_no_twiddle~107_combout ;
wire \reg_no_twiddle[2][1][0]~q ;
wire \reg_no_twiddle~97_combout ;
wire \reg_no_twiddle[3][1][0]~q ;
wire \reg_no_twiddle~87_combout ;
wire \reg_no_twiddle[4][1][0]~q ;
wire \reg_no_twiddle~75_combout ;
wire \reg_no_twiddle[5][1][0]~q ;
wire \reg_no_twiddle~55_combout ;
wire \reg_no_twiddle[0][0][4]~1_combout ;
wire \reg_no_twiddle[0][0][4]~q ;
wire \reg_no_twiddle~118_combout ;
wire \reg_no_twiddle[1][0][4]~q ;
wire \reg_no_twiddle~108_combout ;
wire \reg_no_twiddle[2][0][4]~q ;
wire \reg_no_twiddle~98_combout ;
wire \reg_no_twiddle[3][0][4]~q ;
wire \reg_no_twiddle~88_combout ;
wire \reg_no_twiddle[4][0][4]~q ;
wire \reg_no_twiddle~76_combout ;
wire \reg_no_twiddle[5][0][4]~q ;
wire \reg_no_twiddle~56_combout ;
wire \reg_no_twiddle[0][1][4]~1_combout ;
wire \reg_no_twiddle[0][1][4]~q ;
wire \reg_no_twiddle~119_combout ;
wire \reg_no_twiddle[1][1][4]~q ;
wire \reg_no_twiddle~109_combout ;
wire \reg_no_twiddle[2][1][4]~q ;
wire \reg_no_twiddle~99_combout ;
wire \reg_no_twiddle[3][1][4]~q ;
wire \reg_no_twiddle~89_combout ;
wire \reg_no_twiddle[4][1][4]~q ;
wire \reg_no_twiddle~77_combout ;
wire \reg_no_twiddle[5][1][4]~q ;
wire \reg_no_twiddle~57_combout ;
wire \reg_no_twiddle[0][0][3]~1_combout ;
wire \reg_no_twiddle[0][0][3]~q ;
wire \reg_no_twiddle~120_combout ;
wire \reg_no_twiddle[1][0][3]~q ;
wire \reg_no_twiddle~110_combout ;
wire \reg_no_twiddle[2][0][3]~q ;
wire \reg_no_twiddle~100_combout ;
wire \reg_no_twiddle[3][0][3]~q ;
wire \reg_no_twiddle~90_combout ;
wire \reg_no_twiddle[4][0][3]~q ;
wire \reg_no_twiddle~78_combout ;
wire \reg_no_twiddle[5][0][3]~q ;
wire \reg_no_twiddle~58_combout ;
wire \reg_no_twiddle[0][1][3]~1_combout ;
wire \reg_no_twiddle[0][1][3]~q ;
wire \reg_no_twiddle~121_combout ;
wire \reg_no_twiddle[1][1][3]~q ;
wire \reg_no_twiddle~111_combout ;
wire \reg_no_twiddle[2][1][3]~q ;
wire \reg_no_twiddle~101_combout ;
wire \reg_no_twiddle[3][1][3]~q ;
wire \reg_no_twiddle~91_combout ;
wire \reg_no_twiddle[4][1][3]~q ;
wire \reg_no_twiddle~79_combout ;
wire \reg_no_twiddle[5][1][3]~q ;
wire \reg_no_twiddle~59_combout ;


fftsign_asj_fft_pround_7 \gen_full_rnd:gen_rounding_blk:0:u1 (
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2018(\butterfly_st2[0][1][8]~q ),
	.butterfly_st2017(\butterfly_st2[0][1][7]~q ),
	.butterfly_st2016(\butterfly_st2[0][1][6]~q ),
	.butterfly_st2015(\butterfly_st2[0][1][5]~q ),
	.butterfly_st2014(\butterfly_st2[0][1][4]~q ),
	.butterfly_st2013(\butterfly_st2[0][1][3]~q ),
	.butterfly_st2012(\butterfly_st2[0][1][2]~q ),
	.butterfly_st2011(\butterfly_st2[0][1][1]~q ),
	.butterfly_st2010(\butterfly_st2[0][1][0]~q ),
	.butterfly_st20111(\butterfly_st2[0][1][11]~q ),
	.butterfly_st20110(\butterfly_st2[0][1][10]~q ),
	.butterfly_st2019(\butterfly_st2[0][1][9]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_6 \gen_full_rnd:gen_rounding_blk:0:u0 (
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.butterfly_st2008(\butterfly_st2[0][0][8]~q ),
	.butterfly_st2007(\butterfly_st2[0][0][7]~q ),
	.butterfly_st2006(\butterfly_st2[0][0][6]~q ),
	.butterfly_st2005(\butterfly_st2[0][0][5]~q ),
	.butterfly_st2004(\butterfly_st2[0][0][4]~q ),
	.butterfly_st2003(\butterfly_st2[0][0][3]~q ),
	.butterfly_st2002(\butterfly_st2[0][0][2]~q ),
	.butterfly_st2001(\butterfly_st2[0][0][1]~q ),
	.butterfly_st2000(\butterfly_st2[0][0][0]~q ),
	.butterfly_st20011(\butterfly_st2[0][0][11]~q ),
	.butterfly_st20010(\butterfly_st2[0][0][10]~q ),
	.butterfly_st2009(\butterfly_st2[0][0][9]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_cmult_std_2 \gen_da0:gen_std:cm3 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_14),
	.tdl_arr_9_1(tdl_arr_9_14),
	.tdl_arr_5_11(tdl_arr_5_15),
	.tdl_arr_9_11(tdl_arr_9_15),
	.tdl_arr_6_1(tdl_arr_6_14),
	.tdl_arr_6_11(tdl_arr_6_15),
	.tdl_arr_7_1(tdl_arr_7_14),
	.tdl_arr_7_11(tdl_arr_7_15),
	.tdl_arr_8_1(tdl_arr_8_14),
	.tdl_arr_8_11(tdl_arr_8_15),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_2_11(tdl_arr_2_13),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_1_11(tdl_arr_1_13),
	.tdl_arr_0_1(tdl_arr_0_1),
	.tdl_arr_0_11(tdl_arr_0_13),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_4_11(tdl_arr_4_13),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_3_11(tdl_arr_3_13),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.twiddle_data218(twiddle_data218),
	.twiddle_data219(twiddle_data219),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data208(twiddle_data208),
	.twiddle_data209(twiddle_data209),
	.clk(clk));

fftsign_asj_fft_cmult_std_1 \gen_da0:gen_std:cm2 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_12),
	.tdl_arr_9_1(tdl_arr_9_12),
	.tdl_arr_5_11(tdl_arr_5_13),
	.tdl_arr_9_11(tdl_arr_9_13),
	.tdl_arr_6_1(tdl_arr_6_12),
	.tdl_arr_6_11(tdl_arr_6_13),
	.tdl_arr_7_1(tdl_arr_7_12),
	.tdl_arr_7_11(tdl_arr_7_13),
	.tdl_arr_8_1(tdl_arr_8_12),
	.tdl_arr_8_11(tdl_arr_8_13),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_2_11(tdl_arr_2_14),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_1_11(tdl_arr_1_14),
	.tdl_arr_0_1(tdl_arr_0_11),
	.tdl_arr_0_11(tdl_arr_0_14),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_4_11(tdl_arr_4_14),
	.tdl_arr_3_1(tdl_arr_3_11),
	.tdl_arr_3_11(tdl_arr_3_14),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.twiddle_data118(twiddle_data118),
	.twiddle_data119(twiddle_data119),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data108(twiddle_data108),
	.twiddle_data109(twiddle_data109),
	.clk(clk));

fftsign_asj_fft_cmult_std \gen_da0:gen_std:cm1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_9_1(tdl_arr_9_1),
	.tdl_arr_5_11(tdl_arr_5_11),
	.tdl_arr_9_11(tdl_arr_9_11),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_6_11(tdl_arr_6_11),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_7_11(tdl_arr_7_11),
	.tdl_arr_8_1(tdl_arr_8_1),
	.tdl_arr_8_11(tdl_arr_8_11),
	.tdl_arr_2_1(tdl_arr_2_12),
	.tdl_arr_2_11(tdl_arr_2_15),
	.tdl_arr_1_1(tdl_arr_1_12),
	.tdl_arr_1_11(tdl_arr_1_15),
	.tdl_arr_0_1(tdl_arr_0_12),
	.tdl_arr_0_11(tdl_arr_0_15),
	.tdl_arr_4_1(tdl_arr_4_12),
	.tdl_arr_4_11(tdl_arr_4_15),
	.tdl_arr_3_1(tdl_arr_3_12),
	.tdl_arr_3_11(tdl_arr_3_15),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data018(twiddle_data018),
	.twiddle_data019(twiddle_data019),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data008(twiddle_data008),
	.twiddle_data009(twiddle_data009),
	.clk(clk));

fftsign_asj_fft_bfp_i \gen_disc:bfp_scale (
	.r_array_out_7_2(\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.r_array_out_7_0(\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.r_array_out_6_2(\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.r_array_out_6_0(\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.r_array_out_5_2(\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.r_array_out_5_0(\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.r_array_out_4_2(\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.r_array_out_4_0(\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.r_array_out_3_2(\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.r_array_out_3_0(\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.r_array_out_2_2(\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.r_array_out_2_0(\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.r_array_out_7_3(\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.r_array_out_7_1(\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.r_array_out_6_3(\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.r_array_out_6_1(\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.r_array_out_5_3(\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.r_array_out_5_1(\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.r_array_out_4_3(\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.r_array_out_4_1(\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.r_array_out_3_3(\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.r_array_out_3_1(\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.r_array_out_2_3(\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.r_array_out_2_1(\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.i_array_out_7_2(\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.i_array_out_7_0(\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.i_array_out_6_2(\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.i_array_out_6_0(\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.i_array_out_5_2(\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.i_array_out_5_0(\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.i_array_out_4_2(\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.i_array_out_4_0(\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.i_array_out_3_2(\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.i_array_out_3_0(\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.i_array_out_2_2(\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.i_array_out_2_0(\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.i_array_out_7_3(\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.i_array_out_7_1(\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.i_array_out_6_3(\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.i_array_out_6_1(\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.i_array_out_5_3(\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.i_array_out_5_1(\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.i_array_out_4_3(\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.i_array_out_4_1(\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.i_array_out_3_3(\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.i_array_out_3_1(\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.i_array_out_2_3(\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.i_array_out_2_1(\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_8_0(ram_in_reg_8_0),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_8_2(ram_in_reg_8_2),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_8_1(ram_in_reg_8_1),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_8_3(ram_in_reg_8_3),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_9_0(ram_in_reg_9_0),
	.ram_in_reg_9_2(ram_in_reg_9_2),
	.ram_in_reg_9_1(ram_in_reg_9_1),
	.ram_in_reg_9_3(ram_in_reg_9_3),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_8_4(ram_in_reg_8_4),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_8_6(ram_in_reg_8_6),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_8_5(ram_in_reg_8_5),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_8_7(ram_in_reg_8_7),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.ram_in_reg_9_4(ram_in_reg_9_4),
	.ram_in_reg_9_6(ram_in_reg_9_6),
	.ram_in_reg_9_5(ram_in_reg_9_5),
	.ram_in_reg_9_7(ram_in_reg_9_7),
	.global_clock_enable(global_clock_enable),
	.slb_last_0(slb_last_0),
	.slb_last_1(slb_last_1),
	.slb_last_2(slb_last_2),
	.r_array_out_8_0(\gen_disc:bfp_scale|r_array_out[0][8]~q ),
	.r_array_out_8_2(\gen_disc:bfp_scale|r_array_out[2][8]~q ),
	.r_array_out_1_0(\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.r_array_out_1_2(\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.r_array_out_0_0(\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.r_array_out_0_2(\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.r_array_out_8_1(\gen_disc:bfp_scale|r_array_out[1][8]~q ),
	.r_array_out_8_3(\gen_disc:bfp_scale|r_array_out[3][8]~q ),
	.r_array_out_1_1(\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.r_array_out_1_3(\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.r_array_out_0_1(\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.r_array_out_0_3(\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.r_array_out_9_0(\gen_disc:bfp_scale|r_array_out[0][9]~q ),
	.r_array_out_9_2(\gen_disc:bfp_scale|r_array_out[2][9]~q ),
	.r_array_out_9_1(\gen_disc:bfp_scale|r_array_out[1][9]~q ),
	.r_array_out_9_3(\gen_disc:bfp_scale|r_array_out[3][9]~q ),
	.i_array_out_8_0(\gen_disc:bfp_scale|i_array_out[0][8]~q ),
	.i_array_out_8_2(\gen_disc:bfp_scale|i_array_out[2][8]~q ),
	.i_array_out_1_0(\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.i_array_out_1_2(\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.i_array_out_0_0(\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.i_array_out_0_2(\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.i_array_out_8_1(\gen_disc:bfp_scale|i_array_out[1][8]~q ),
	.i_array_out_8_3(\gen_disc:bfp_scale|i_array_out[3][8]~q ),
	.i_array_out_1_1(\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.i_array_out_1_3(\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.i_array_out_0_1(\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.i_array_out_0_3(\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.i_array_out_9_0(\gen_disc:bfp_scale|i_array_out[0][9]~q ),
	.i_array_out_9_2(\gen_disc:bfp_scale|i_array_out[2][9]~q ),
	.i_array_out_9_1(\gen_disc:bfp_scale|i_array_out[1][9]~q ),
	.i_array_out_9_3(\gen_disc:bfp_scale|i_array_out[3][9]~q ),
	.clk(clk));

fftsign_asj_fft_bfp_o \gen_disc:bfp_detect (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(tdl_arr_0),
	.sdetdIDLE(sdetdIDLE),
	.slb_i_0(slb_i_0),
	.slb_i_1(slb_i_1),
	.slb_i_2(slb_i_2),
	.slb_i_3(slb_i_3),
	.Mux2(Mux2),
	.Mux1(Mux1),
	.tdl_arr_6(tdl_arr_6),
	.reg_no_twiddle605(reg_no_twiddle605),
	.reg_no_twiddle609(reg_no_twiddle609),
	.reg_no_twiddle615(reg_no_twiddle615),
	.reg_no_twiddle619(reg_no_twiddle619),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_9_1(tdl_arr_9_1),
	.tdl_arr_5_11(tdl_arr_5_11),
	.tdl_arr_9_11(tdl_arr_9_11),
	.tdl_arr_5_12(tdl_arr_5_12),
	.tdl_arr_9_12(tdl_arr_9_12),
	.tdl_arr_5_13(tdl_arr_5_13),
	.tdl_arr_9_13(tdl_arr_9_13),
	.tdl_arr_5_14(tdl_arr_5_14),
	.tdl_arr_9_14(tdl_arr_9_14),
	.tdl_arr_5_15(tdl_arr_5_15),
	.tdl_arr_9_15(tdl_arr_9_15),
	.reg_no_twiddle606(reg_no_twiddle606),
	.reg_no_twiddle616(reg_no_twiddle616),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_6_11(tdl_arr_6_11),
	.tdl_arr_6_12(tdl_arr_6_12),
	.tdl_arr_6_13(tdl_arr_6_13),
	.tdl_arr_6_14(tdl_arr_6_14),
	.tdl_arr_6_15(tdl_arr_6_15),
	.reg_no_twiddle607(reg_no_twiddle607),
	.reg_no_twiddle617(reg_no_twiddle617),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_7_11(tdl_arr_7_11),
	.tdl_arr_7_12(tdl_arr_7_12),
	.tdl_arr_7_13(tdl_arr_7_13),
	.tdl_arr_7_14(tdl_arr_7_14),
	.tdl_arr_7_15(tdl_arr_7_15),
	.reg_no_twiddle608(reg_no_twiddle608),
	.reg_no_twiddle618(reg_no_twiddle618),
	.tdl_arr_8_1(tdl_arr_8_1),
	.tdl_arr_8_11(tdl_arr_8_11),
	.tdl_arr_8_12(tdl_arr_8_12),
	.tdl_arr_8_13(tdl_arr_8_13),
	.tdl_arr_8_14(tdl_arr_8_14),
	.tdl_arr_8_15(tdl_arr_8_15),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_pround_13 \gen_full_rnd:gen_rounding_blk:3:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2312(\butterfly_st2[3][1][2]~q ),
	.butterfly_st2311(\butterfly_st2[3][1][1]~q ),
	.butterfly_st2310(\butterfly_st2[3][1][0]~q ),
	.butterfly_st23111(\butterfly_st2[3][1][11]~q ),
	.butterfly_st2313(\butterfly_st2[3][1][3]~q ),
	.butterfly_st2314(\butterfly_st2[3][1][4]~q ),
	.butterfly_st2315(\butterfly_st2[3][1][5]~q ),
	.butterfly_st2316(\butterfly_st2[3][1][6]~q ),
	.butterfly_st2317(\butterfly_st2[3][1][7]~q ),
	.butterfly_st2318(\butterfly_st2[3][1][8]~q ),
	.butterfly_st2319(\butterfly_st2[3][1][9]~q ),
	.butterfly_st23110(\butterfly_st2[3][1][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_12 \gen_full_rnd:gen_rounding_blk:3:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2302(\butterfly_st2[3][0][2]~q ),
	.butterfly_st2301(\butterfly_st2[3][0][1]~q ),
	.butterfly_st2300(\butterfly_st2[3][0][0]~q ),
	.butterfly_st23011(\butterfly_st2[3][0][11]~q ),
	.butterfly_st2303(\butterfly_st2[3][0][3]~q ),
	.butterfly_st2304(\butterfly_st2[3][0][4]~q ),
	.butterfly_st2305(\butterfly_st2[3][0][5]~q ),
	.butterfly_st2306(\butterfly_st2[3][0][6]~q ),
	.butterfly_st2307(\butterfly_st2[3][0][7]~q ),
	.butterfly_st2308(\butterfly_st2[3][0][8]~q ),
	.butterfly_st2309(\butterfly_st2[3][0][9]~q ),
	.butterfly_st23010(\butterfly_st2[3][0][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_11 \gen_full_rnd:gen_rounding_blk:2:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2212(\butterfly_st2[2][1][2]~q ),
	.butterfly_st2211(\butterfly_st2[2][1][1]~q ),
	.butterfly_st2210(\butterfly_st2[2][1][0]~q ),
	.butterfly_st22111(\butterfly_st2[2][1][11]~q ),
	.butterfly_st2213(\butterfly_st2[2][1][3]~q ),
	.butterfly_st2214(\butterfly_st2[2][1][4]~q ),
	.butterfly_st2215(\butterfly_st2[2][1][5]~q ),
	.butterfly_st2216(\butterfly_st2[2][1][6]~q ),
	.butterfly_st2217(\butterfly_st2[2][1][7]~q ),
	.butterfly_st2218(\butterfly_st2[2][1][8]~q ),
	.butterfly_st2219(\butterfly_st2[2][1][9]~q ),
	.butterfly_st22110(\butterfly_st2[2][1][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_10 \gen_full_rnd:gen_rounding_blk:2:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2202(\butterfly_st2[2][0][2]~q ),
	.butterfly_st2201(\butterfly_st2[2][0][1]~q ),
	.butterfly_st2200(\butterfly_st2[2][0][0]~q ),
	.butterfly_st22011(\butterfly_st2[2][0][11]~q ),
	.butterfly_st2203(\butterfly_st2[2][0][3]~q ),
	.butterfly_st2204(\butterfly_st2[2][0][4]~q ),
	.butterfly_st2205(\butterfly_st2[2][0][5]~q ),
	.butterfly_st2206(\butterfly_st2[2][0][6]~q ),
	.butterfly_st2207(\butterfly_st2[2][0][7]~q ),
	.butterfly_st2208(\butterfly_st2[2][0][8]~q ),
	.butterfly_st2209(\butterfly_st2[2][0][9]~q ),
	.butterfly_st22010(\butterfly_st2[2][0][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_9 \gen_full_rnd:gen_rounding_blk:1:u1 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2112(\butterfly_st2[1][1][2]~q ),
	.butterfly_st2111(\butterfly_st2[1][1][1]~q ),
	.butterfly_st2110(\butterfly_st2[1][1][0]~q ),
	.butterfly_st21111(\butterfly_st2[1][1][11]~q ),
	.butterfly_st2113(\butterfly_st2[1][1][3]~q ),
	.butterfly_st2114(\butterfly_st2[1][1][4]~q ),
	.butterfly_st2115(\butterfly_st2[1][1][5]~q ),
	.butterfly_st2116(\butterfly_st2[1][1][6]~q ),
	.butterfly_st2117(\butterfly_st2[1][1][7]~q ),
	.butterfly_st2118(\butterfly_st2[1][1][8]~q ),
	.butterfly_st2119(\butterfly_st2[1][1][9]~q ),
	.butterfly_st21110(\butterfly_st2[1][1][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_8 \gen_full_rnd:gen_rounding_blk:1:u0 (
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.butterfly_st2102(\butterfly_st2[1][0][2]~q ),
	.butterfly_st2101(\butterfly_st2[1][0][1]~q ),
	.butterfly_st2100(\butterfly_st2[1][0][0]~q ),
	.butterfly_st21011(\butterfly_st2[1][0][11]~q ),
	.butterfly_st2103(\butterfly_st2[1][0][3]~q ),
	.butterfly_st2104(\butterfly_st2[1][0][4]~q ),
	.butterfly_st2105(\butterfly_st2[1][0][5]~q ),
	.butterfly_st2106(\butterfly_st2[1][0][6]~q ),
	.butterfly_st2107(\butterfly_st2[1][0][7]~q ),
	.butterfly_st2108(\butterfly_st2[1][0][8]~q ),
	.butterfly_st2109(\butterfly_st2[1][0][9]~q ),
	.butterfly_st21010(\butterfly_st2[1][0][10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

dffeas \butterfly_st2[0][0][8] (
	.clk(clk),
	.d(\butterfly_st2[0][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][8] .power_up = "low";

dffeas \butterfly_st2[0][0][7] (
	.clk(clk),
	.d(\butterfly_st2[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][7] .power_up = "low";

dffeas \butterfly_st2[0][0][6] (
	.clk(clk),
	.d(\butterfly_st2[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][6] .power_up = "low";

dffeas \butterfly_st2[0][0][5] (
	.clk(clk),
	.d(\butterfly_st2[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][5] .power_up = "low";

dffeas \butterfly_st2[0][0][4] (
	.clk(clk),
	.d(\butterfly_st2[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][4] .power_up = "low";

dffeas \butterfly_st2[0][0][3] (
	.clk(clk),
	.d(\butterfly_st2[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][3] .power_up = "low";

dffeas \butterfly_st2[0][0][2] (
	.clk(clk),
	.d(\butterfly_st2[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][2] .power_up = "low";

dffeas \butterfly_st2[0][0][1] (
	.clk(clk),
	.d(\butterfly_st2[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][1] .power_up = "low";

dffeas \butterfly_st2[0][0][0] (
	.clk(clk),
	.d(\butterfly_st2[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][0] .power_up = "low";

dffeas \butterfly_st2[0][0][11] (
	.clk(clk),
	.d(\butterfly_st2[0][0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][11] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][11] .power_up = "low";

dffeas \butterfly_st2[0][0][10] (
	.clk(clk),
	.d(\butterfly_st2[0][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][10] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][10] .power_up = "low";

dffeas \butterfly_st2[0][0][9] (
	.clk(clk),
	.d(\butterfly_st2[0][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][9] .power_up = "low";

dffeas \butterfly_st2[0][1][8] (
	.clk(clk),
	.d(\butterfly_st2[0][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][8] .power_up = "low";

dffeas \butterfly_st2[0][1][7] (
	.clk(clk),
	.d(\butterfly_st2[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][7] .power_up = "low";

dffeas \butterfly_st2[0][1][6] (
	.clk(clk),
	.d(\butterfly_st2[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][6] .power_up = "low";

dffeas \butterfly_st2[0][1][5] (
	.clk(clk),
	.d(\butterfly_st2[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][5] .power_up = "low";

dffeas \butterfly_st2[0][1][4] (
	.clk(clk),
	.d(\butterfly_st2[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][4] .power_up = "low";

dffeas \butterfly_st2[0][1][3] (
	.clk(clk),
	.d(\butterfly_st2[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][3] .power_up = "low";

dffeas \butterfly_st2[0][1][2] (
	.clk(clk),
	.d(\butterfly_st2[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][2] .power_up = "low";

dffeas \butterfly_st2[0][1][1] (
	.clk(clk),
	.d(\butterfly_st2[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][1] .power_up = "low";

dffeas \butterfly_st2[0][1][0] (
	.clk(clk),
	.d(\butterfly_st2[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][0] .power_up = "low";

dffeas \butterfly_st2[0][1][11] (
	.clk(clk),
	.d(\butterfly_st2[0][1][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][11] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][11] .power_up = "low";

dffeas \butterfly_st2[0][1][10] (
	.clk(clk),
	.d(\butterfly_st2[0][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][10] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][10] .power_up = "low";

dffeas \butterfly_st2[0][1][9] (
	.clk(clk),
	.d(\butterfly_st2[0][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[0][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][9] .power_up = "low";

dffeas \butterfly_st2[1][1][2] (
	.clk(clk),
	.d(\butterfly_st2[1][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][2] .power_up = "low";

dffeas \butterfly_st2[1][1][1] (
	.clk(clk),
	.d(\butterfly_st2[1][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][1] .power_up = "low";

dffeas \butterfly_st2[1][1][0] (
	.clk(clk),
	.d(\butterfly_st2[1][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][0] .power_up = "low";

dffeas \butterfly_st2[1][1][11] (
	.clk(clk),
	.d(\butterfly_st2[1][1][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][11] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][11] .power_up = "low";

dffeas \butterfly_st2[1][1][3] (
	.clk(clk),
	.d(\butterfly_st2[1][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][3] .power_up = "low";

dffeas \butterfly_st2[1][1][4] (
	.clk(clk),
	.d(\butterfly_st2[1][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][4] .power_up = "low";

dffeas \butterfly_st2[1][1][5] (
	.clk(clk),
	.d(\butterfly_st2[1][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][5] .power_up = "low";

dffeas \butterfly_st2[1][1][6] (
	.clk(clk),
	.d(\butterfly_st2[1][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][6] .power_up = "low";

dffeas \butterfly_st2[1][1][7] (
	.clk(clk),
	.d(\butterfly_st2[1][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][7] .power_up = "low";

dffeas \butterfly_st2[1][1][8] (
	.clk(clk),
	.d(\butterfly_st2[1][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][8] .power_up = "low";

dffeas \butterfly_st2[1][1][9] (
	.clk(clk),
	.d(\butterfly_st2[1][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][9] .power_up = "low";

dffeas \butterfly_st2[1][1][10] (
	.clk(clk),
	.d(\butterfly_st2[1][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][10] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][10] .power_up = "low";

dffeas \butterfly_st2[1][0][2] (
	.clk(clk),
	.d(\butterfly_st2[1][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][2] .power_up = "low";

dffeas \butterfly_st2[1][0][1] (
	.clk(clk),
	.d(\butterfly_st2[1][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][1] .power_up = "low";

dffeas \butterfly_st2[1][0][0] (
	.clk(clk),
	.d(\butterfly_st2[1][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][0] .power_up = "low";

dffeas \butterfly_st2[1][0][11] (
	.clk(clk),
	.d(\butterfly_st2[1][0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][11] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][11] .power_up = "low";

dffeas \butterfly_st2[1][0][3] (
	.clk(clk),
	.d(\butterfly_st2[1][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][3] .power_up = "low";

dffeas \butterfly_st2[1][0][4] (
	.clk(clk),
	.d(\butterfly_st2[1][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][4] .power_up = "low";

dffeas \butterfly_st2[1][0][5] (
	.clk(clk),
	.d(\butterfly_st2[1][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][5] .power_up = "low";

dffeas \butterfly_st2[1][0][6] (
	.clk(clk),
	.d(\butterfly_st2[1][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][6] .power_up = "low";

dffeas \butterfly_st2[1][0][7] (
	.clk(clk),
	.d(\butterfly_st2[1][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][7] .power_up = "low";

dffeas \butterfly_st2[1][0][8] (
	.clk(clk),
	.d(\butterfly_st2[1][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][8] .power_up = "low";

dffeas \butterfly_st2[1][0][9] (
	.clk(clk),
	.d(\butterfly_st2[1][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][9] .power_up = "low";

dffeas \butterfly_st2[1][0][10] (
	.clk(clk),
	.d(\butterfly_st2[1][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[1][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][10] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][10] .power_up = "low";

dffeas \butterfly_st2[2][1][2] (
	.clk(clk),
	.d(\butterfly_st2[2][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][2] .power_up = "low";

dffeas \butterfly_st2[2][1][1] (
	.clk(clk),
	.d(\butterfly_st2[2][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][1] .power_up = "low";

dffeas \butterfly_st2[2][1][0] (
	.clk(clk),
	.d(\butterfly_st2[2][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][0] .power_up = "low";

dffeas \butterfly_st2[2][1][11] (
	.clk(clk),
	.d(\butterfly_st2[2][1][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][11] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][11] .power_up = "low";

dffeas \butterfly_st2[2][1][3] (
	.clk(clk),
	.d(\butterfly_st2[2][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][3] .power_up = "low";

dffeas \butterfly_st2[2][1][4] (
	.clk(clk),
	.d(\butterfly_st2[2][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][4] .power_up = "low";

dffeas \butterfly_st2[2][1][5] (
	.clk(clk),
	.d(\butterfly_st2[2][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][5] .power_up = "low";

dffeas \butterfly_st2[2][1][6] (
	.clk(clk),
	.d(\butterfly_st2[2][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][6] .power_up = "low";

dffeas \butterfly_st2[2][1][7] (
	.clk(clk),
	.d(\butterfly_st2[2][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][7] .power_up = "low";

dffeas \butterfly_st2[2][1][8] (
	.clk(clk),
	.d(\butterfly_st2[2][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][8] .power_up = "low";

dffeas \butterfly_st2[2][1][9] (
	.clk(clk),
	.d(\butterfly_st2[2][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][9] .power_up = "low";

dffeas \butterfly_st2[2][1][10] (
	.clk(clk),
	.d(\butterfly_st2[2][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][10] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][10] .power_up = "low";

dffeas \butterfly_st2[2][0][2] (
	.clk(clk),
	.d(\butterfly_st2[2][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][2] .power_up = "low";

dffeas \butterfly_st2[2][0][1] (
	.clk(clk),
	.d(\butterfly_st2[2][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][1] .power_up = "low";

dffeas \butterfly_st2[2][0][0] (
	.clk(clk),
	.d(\butterfly_st2[2][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][0] .power_up = "low";

dffeas \butterfly_st2[2][0][11] (
	.clk(clk),
	.d(\butterfly_st2[2][0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][11] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][11] .power_up = "low";

dffeas \butterfly_st2[2][0][3] (
	.clk(clk),
	.d(\butterfly_st2[2][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][3] .power_up = "low";

dffeas \butterfly_st2[2][0][4] (
	.clk(clk),
	.d(\butterfly_st2[2][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][4] .power_up = "low";

dffeas \butterfly_st2[2][0][5] (
	.clk(clk),
	.d(\butterfly_st2[2][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][5] .power_up = "low";

dffeas \butterfly_st2[2][0][6] (
	.clk(clk),
	.d(\butterfly_st2[2][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][6] .power_up = "low";

dffeas \butterfly_st2[2][0][7] (
	.clk(clk),
	.d(\butterfly_st2[2][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][7] .power_up = "low";

dffeas \butterfly_st2[2][0][8] (
	.clk(clk),
	.d(\butterfly_st2[2][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][8] .power_up = "low";

dffeas \butterfly_st2[2][0][9] (
	.clk(clk),
	.d(\butterfly_st2[2][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][9] .power_up = "low";

dffeas \butterfly_st2[2][0][10] (
	.clk(clk),
	.d(\butterfly_st2[2][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[2][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][10] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][10] .power_up = "low";

dffeas \butterfly_st2[3][1][2] (
	.clk(clk),
	.d(\butterfly_st2[3][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][2] .power_up = "low";

dffeas \butterfly_st2[3][1][1] (
	.clk(clk),
	.d(\butterfly_st2[3][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][1] .power_up = "low";

dffeas \butterfly_st2[3][1][0] (
	.clk(clk),
	.d(\butterfly_st2[3][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][0] .power_up = "low";

dffeas \butterfly_st2[3][1][11] (
	.clk(clk),
	.d(\butterfly_st2[3][1][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][11] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][11] .power_up = "low";

dffeas \butterfly_st2[3][1][3] (
	.clk(clk),
	.d(\butterfly_st2[3][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][3] .power_up = "low";

dffeas \butterfly_st2[3][1][4] (
	.clk(clk),
	.d(\butterfly_st2[3][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][4] .power_up = "low";

dffeas \butterfly_st2[3][1][5] (
	.clk(clk),
	.d(\butterfly_st2[3][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][5] .power_up = "low";

dffeas \butterfly_st2[3][1][6] (
	.clk(clk),
	.d(\butterfly_st2[3][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][6] .power_up = "low";

dffeas \butterfly_st2[3][1][7] (
	.clk(clk),
	.d(\butterfly_st2[3][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][7] .power_up = "low";

dffeas \butterfly_st2[3][1][8] (
	.clk(clk),
	.d(\butterfly_st2[3][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][8] .power_up = "low";

dffeas \butterfly_st2[3][1][9] (
	.clk(clk),
	.d(\butterfly_st2[3][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][9] .power_up = "low";

dffeas \butterfly_st2[3][1][10] (
	.clk(clk),
	.d(\butterfly_st2[3][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][10] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][10] .power_up = "low";

dffeas \butterfly_st2[3][0][2] (
	.clk(clk),
	.d(\butterfly_st2[3][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][2] .power_up = "low";

dffeas \butterfly_st2[3][0][1] (
	.clk(clk),
	.d(\butterfly_st2[3][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][1] .power_up = "low";

dffeas \butterfly_st2[3][0][0] (
	.clk(clk),
	.d(\butterfly_st2[3][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][0] .power_up = "low";

dffeas \butterfly_st2[3][0][11] (
	.clk(clk),
	.d(\butterfly_st2[3][0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][11]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][11] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][11] .power_up = "low";

dffeas \butterfly_st2[3][0][3] (
	.clk(clk),
	.d(\butterfly_st2[3][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][3] .power_up = "low";

dffeas \butterfly_st2[3][0][4] (
	.clk(clk),
	.d(\butterfly_st2[3][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][4] .power_up = "low";

dffeas \butterfly_st2[3][0][5] (
	.clk(clk),
	.d(\butterfly_st2[3][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][5] .power_up = "low";

dffeas \butterfly_st2[3][0][6] (
	.clk(clk),
	.d(\butterfly_st2[3][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][6] .power_up = "low";

dffeas \butterfly_st2[3][0][7] (
	.clk(clk),
	.d(\butterfly_st2[3][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][7] .power_up = "low";

dffeas \butterfly_st2[3][0][8] (
	.clk(clk),
	.d(\butterfly_st2[3][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][8] .power_up = "low";

dffeas \butterfly_st2[3][0][9] (
	.clk(clk),
	.d(\butterfly_st2[3][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][9] .power_up = "low";

dffeas \butterfly_st2[3][0][10] (
	.clk(clk),
	.d(\butterfly_st2[3][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st2[3][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][10] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][10] .power_up = "low";

dffeas \butterfly_st1[0][0][8] (
	.clk(clk),
	.d(\butterfly_st1[0][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][8] .power_up = "low";

dffeas \butterfly_st1[1][0][8] (
	.clk(clk),
	.d(\butterfly_st1[1][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][7] (
	.clk(clk),
	.d(\butterfly_st1[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][7] .power_up = "low";

dffeas \butterfly_st1[1][0][7] (
	.clk(clk),
	.d(\butterfly_st1[1][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][7] .power_up = "low";

dffeas \butterfly_st1[0][0][6] (
	.clk(clk),
	.d(\butterfly_st1[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][6] .power_up = "low";

dffeas \butterfly_st1[1][0][6] (
	.clk(clk),
	.d(\butterfly_st1[1][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][6] .power_up = "low";

dffeas \butterfly_st1[0][0][5] (
	.clk(clk),
	.d(\butterfly_st1[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][5] .power_up = "low";

dffeas \butterfly_st1[1][0][5] (
	.clk(clk),
	.d(\butterfly_st1[1][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][5] .power_up = "low";

dffeas \butterfly_st1[0][0][4] (
	.clk(clk),
	.d(\butterfly_st1[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][4] .power_up = "low";

dffeas \butterfly_st1[1][0][4] (
	.clk(clk),
	.d(\butterfly_st1[1][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][4] .power_up = "low";

dffeas \butterfly_st1[0][0][3] (
	.clk(clk),
	.d(\butterfly_st1[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][3] .power_up = "low";

dffeas \butterfly_st1[1][0][3] (
	.clk(clk),
	.d(\butterfly_st1[1][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][3] .power_up = "low";

dffeas \butterfly_st1[0][0][2] (
	.clk(clk),
	.d(\butterfly_st1[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][2] .power_up = "low";

dffeas \butterfly_st1[1][0][2] (
	.clk(clk),
	.d(\butterfly_st1[1][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][2] .power_up = "low";

dffeas \butterfly_st1[0][0][1] (
	.clk(clk),
	.d(\butterfly_st1[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][1] .power_up = "low";

dffeas \butterfly_st1[1][0][1] (
	.clk(clk),
	.d(\butterfly_st1[1][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][1] .power_up = "low";

dffeas \butterfly_st1[0][0][0] (
	.clk(clk),
	.d(\butterfly_st1[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][0] .power_up = "low";

dffeas \butterfly_st1[1][0][0] (
	.clk(clk),
	.d(\butterfly_st1[1][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[0][0][0]~1 (
	.dataa(\butterfly_st1[0][0][0]~q ),
	.datab(\butterfly_st1[1][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[0][0][0]~1_combout ),
	.cout(\butterfly_st2[0][0][0]~2 ));
defparam \butterfly_st2[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[0][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[0][0][1]~1 (
	.dataa(\butterfly_st1[0][0][1]~q ),
	.datab(\butterfly_st1[1][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][0]~2 ),
	.combout(\butterfly_st2[0][0][1]~1_combout ),
	.cout(\butterfly_st2[0][0][1]~2 ));
defparam \butterfly_st2[0][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][2]~1 (
	.dataa(\butterfly_st1[0][0][2]~q ),
	.datab(\butterfly_st1[1][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][1]~2 ),
	.combout(\butterfly_st2[0][0][2]~1_combout ),
	.cout(\butterfly_st2[0][0][2]~2 ));
defparam \butterfly_st2[0][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][3]~1 (
	.dataa(\butterfly_st1[0][0][3]~q ),
	.datab(\butterfly_st1[1][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][2]~2 ),
	.combout(\butterfly_st2[0][0][3]~1_combout ),
	.cout(\butterfly_st2[0][0][3]~2 ));
defparam \butterfly_st2[0][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][4]~1 (
	.dataa(\butterfly_st1[0][0][4]~q ),
	.datab(\butterfly_st1[1][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][3]~2 ),
	.combout(\butterfly_st2[0][0][4]~1_combout ),
	.cout(\butterfly_st2[0][0][4]~2 ));
defparam \butterfly_st2[0][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][5]~1 (
	.dataa(\butterfly_st1[0][0][5]~q ),
	.datab(\butterfly_st1[1][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][4]~2 ),
	.combout(\butterfly_st2[0][0][5]~1_combout ),
	.cout(\butterfly_st2[0][0][5]~2 ));
defparam \butterfly_st2[0][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][6]~1 (
	.dataa(\butterfly_st1[0][0][6]~q ),
	.datab(\butterfly_st1[1][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][5]~2 ),
	.combout(\butterfly_st2[0][0][6]~1_combout ),
	.cout(\butterfly_st2[0][0][6]~2 ));
defparam \butterfly_st2[0][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][7]~1 (
	.dataa(\butterfly_st1[0][0][7]~q ),
	.datab(\butterfly_st1[1][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][6]~2 ),
	.combout(\butterfly_st2[0][0][7]~1_combout ),
	.cout(\butterfly_st2[0][0][7]~2 ));
defparam \butterfly_st2[0][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][8]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][7]~2 ),
	.combout(\butterfly_st2[0][0][8]~1_combout ),
	.cout(\butterfly_st2[0][0][8]~2 ));
defparam \butterfly_st2[0][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][8]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[0][0][10] (
	.clk(clk),
	.d(\butterfly_st1[0][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][10] .power_up = "low";

dffeas \butterfly_st1[1][0][10] (
	.clk(clk),
	.d(\butterfly_st1[1][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][10] .power_up = "low";

dffeas \butterfly_st1[0][0][9] (
	.clk(clk),
	.d(\butterfly_st1[0][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][9] .power_up = "low";

dffeas \butterfly_st1[1][0][9] (
	.clk(clk),
	.d(\butterfly_st1[1][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][9] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[0][0][9]~1 (
	.dataa(\butterfly_st1[0][0][9]~q ),
	.datab(\butterfly_st1[1][0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][8]~2 ),
	.combout(\butterfly_st2[0][0][9]~1_combout ),
	.cout(\butterfly_st2[0][0][9]~2 ));
defparam \butterfly_st2[0][0][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][10]~1 (
	.dataa(\butterfly_st1[0][0][10]~q ),
	.datab(\butterfly_st1[1][0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][0][9]~2 ),
	.combout(\butterfly_st2[0][0][10]~1_combout ),
	.cout(\butterfly_st2[0][0][10]~2 ));
defparam \butterfly_st2[0][0][10]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][0][11]~1 (
	.dataa(\butterfly_st1[0][0][10]~q ),
	.datab(\butterfly_st1[1][0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[0][0][10]~2 ),
	.combout(\butterfly_st2[0][0][11]~1_combout ),
	.cout());
defparam \butterfly_st2[0][0][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[0][0][11]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[0][1][8] (
	.clk(clk),
	.d(\butterfly_st1[0][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][8] .power_up = "low";

dffeas \butterfly_st1[1][1][8] (
	.clk(clk),
	.d(\butterfly_st1[1][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][8] .power_up = "low";

dffeas \butterfly_st1[0][1][7] (
	.clk(clk),
	.d(\butterfly_st1[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][7] .power_up = "low";

dffeas \butterfly_st1[1][1][7] (
	.clk(clk),
	.d(\butterfly_st1[1][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][7] .power_up = "low";

dffeas \butterfly_st1[0][1][6] (
	.clk(clk),
	.d(\butterfly_st1[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][6] .power_up = "low";

dffeas \butterfly_st1[1][1][6] (
	.clk(clk),
	.d(\butterfly_st1[1][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][6] .power_up = "low";

dffeas \butterfly_st1[0][1][5] (
	.clk(clk),
	.d(\butterfly_st1[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][5] .power_up = "low";

dffeas \butterfly_st1[1][1][5] (
	.clk(clk),
	.d(\butterfly_st1[1][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][5] .power_up = "low";

dffeas \butterfly_st1[0][1][4] (
	.clk(clk),
	.d(\butterfly_st1[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][4] .power_up = "low";

dffeas \butterfly_st1[1][1][4] (
	.clk(clk),
	.d(\butterfly_st1[1][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][4] .power_up = "low";

dffeas \butterfly_st1[0][1][3] (
	.clk(clk),
	.d(\butterfly_st1[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][3] .power_up = "low";

dffeas \butterfly_st1[1][1][3] (
	.clk(clk),
	.d(\butterfly_st1[1][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][3] .power_up = "low";

dffeas \butterfly_st1[0][1][2] (
	.clk(clk),
	.d(\butterfly_st1[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][2] .power_up = "low";

dffeas \butterfly_st1[1][1][2] (
	.clk(clk),
	.d(\butterfly_st1[1][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][2] .power_up = "low";

dffeas \butterfly_st1[0][1][1] (
	.clk(clk),
	.d(\butterfly_st1[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][1] .power_up = "low";

dffeas \butterfly_st1[1][1][1] (
	.clk(clk),
	.d(\butterfly_st1[1][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][1] .power_up = "low";

dffeas \butterfly_st1[0][1][0] (
	.clk(clk),
	.d(\butterfly_st1[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][0] .power_up = "low";

dffeas \butterfly_st1[1][1][0] (
	.clk(clk),
	.d(\butterfly_st1[1][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[0][1][0]~1 (
	.dataa(\butterfly_st1[0][1][0]~q ),
	.datab(\butterfly_st1[1][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[0][1][0]~1_combout ),
	.cout(\butterfly_st2[0][1][0]~2 ));
defparam \butterfly_st2[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[0][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[0][1][1]~1 (
	.dataa(\butterfly_st1[0][1][1]~q ),
	.datab(\butterfly_st1[1][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][0]~2 ),
	.combout(\butterfly_st2[0][1][1]~1_combout ),
	.cout(\butterfly_st2[0][1][1]~2 ));
defparam \butterfly_st2[0][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][2]~1 (
	.dataa(\butterfly_st1[0][1][2]~q ),
	.datab(\butterfly_st1[1][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][1]~2 ),
	.combout(\butterfly_st2[0][1][2]~1_combout ),
	.cout(\butterfly_st2[0][1][2]~2 ));
defparam \butterfly_st2[0][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][3]~1 (
	.dataa(\butterfly_st1[0][1][3]~q ),
	.datab(\butterfly_st1[1][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][2]~2 ),
	.combout(\butterfly_st2[0][1][3]~1_combout ),
	.cout(\butterfly_st2[0][1][3]~2 ));
defparam \butterfly_st2[0][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][4]~1 (
	.dataa(\butterfly_st1[0][1][4]~q ),
	.datab(\butterfly_st1[1][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][3]~2 ),
	.combout(\butterfly_st2[0][1][4]~1_combout ),
	.cout(\butterfly_st2[0][1][4]~2 ));
defparam \butterfly_st2[0][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][5]~1 (
	.dataa(\butterfly_st1[0][1][5]~q ),
	.datab(\butterfly_st1[1][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][4]~2 ),
	.combout(\butterfly_st2[0][1][5]~1_combout ),
	.cout(\butterfly_st2[0][1][5]~2 ));
defparam \butterfly_st2[0][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][6]~1 (
	.dataa(\butterfly_st1[0][1][6]~q ),
	.datab(\butterfly_st1[1][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][5]~2 ),
	.combout(\butterfly_st2[0][1][6]~1_combout ),
	.cout(\butterfly_st2[0][1][6]~2 ));
defparam \butterfly_st2[0][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][7]~1 (
	.dataa(\butterfly_st1[0][1][7]~q ),
	.datab(\butterfly_st1[1][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][6]~2 ),
	.combout(\butterfly_st2[0][1][7]~1_combout ),
	.cout(\butterfly_st2[0][1][7]~2 ));
defparam \butterfly_st2[0][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][8]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][7]~2 ),
	.combout(\butterfly_st2[0][1][8]~1_combout ),
	.cout(\butterfly_st2[0][1][8]~2 ));
defparam \butterfly_st2[0][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][8]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[0][1][10] (
	.clk(clk),
	.d(\butterfly_st1[0][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][10] .power_up = "low";

dffeas \butterfly_st1[1][1][10] (
	.clk(clk),
	.d(\butterfly_st1[1][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][10] .power_up = "low";

dffeas \butterfly_st1[0][1][9] (
	.clk(clk),
	.d(\butterfly_st1[0][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[0][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][9] .power_up = "low";

dffeas \butterfly_st1[1][1][9] (
	.clk(clk),
	.d(\butterfly_st1[1][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[1][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][9] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[0][1][9]~1 (
	.dataa(\butterfly_st1[0][1][9]~q ),
	.datab(\butterfly_st1[1][1][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][8]~2 ),
	.combout(\butterfly_st2[0][1][9]~1_combout ),
	.cout(\butterfly_st2[0][1][9]~2 ));
defparam \butterfly_st2[0][1][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[0][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][10]~1 (
	.dataa(\butterfly_st1[0][1][10]~q ),
	.datab(\butterfly_st1[1][1][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[0][1][9]~2 ),
	.combout(\butterfly_st2[0][1][10]~1_combout ),
	.cout(\butterfly_st2[0][1][10]~2 ));
defparam \butterfly_st2[0][1][10]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[0][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[0][1][11]~1 (
	.dataa(\butterfly_st1[0][1][10]~q ),
	.datab(\butterfly_st1[1][1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[0][1][10]~2 ),
	.combout(\butterfly_st2[0][1][11]~1_combout ),
	.cout());
defparam \butterfly_st2[0][1][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[0][1][11]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][1][2] (
	.clk(clk),
	.d(\butterfly_st1[2][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][2] .power_up = "low";

dffeas \butterfly_st1[3][0][2] (
	.clk(clk),
	.d(\butterfly_st1[3][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][2] .power_up = "low";

dffeas \butterfly_st1[2][1][1] (
	.clk(clk),
	.d(\butterfly_st1[2][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][1] .power_up = "low";

dffeas \butterfly_st1[3][0][1] (
	.clk(clk),
	.d(\butterfly_st1[3][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][1] .power_up = "low";

dffeas \butterfly_st1[2][1][0] (
	.clk(clk),
	.d(\butterfly_st1[2][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][0] .power_up = "low";

dffeas \butterfly_st1[3][0][0] (
	.clk(clk),
	.d(\butterfly_st1[3][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[1][1][0]~1 (
	.dataa(\butterfly_st1[2][1][0]~q ),
	.datab(\butterfly_st1[3][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[1][1][0]~1_combout ),
	.cout(\butterfly_st2[1][1][0]~2 ));
defparam \butterfly_st2[1][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[1][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[1][1][1]~1 (
	.dataa(\butterfly_st1[2][1][1]~q ),
	.datab(\butterfly_st1[3][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][0]~2 ),
	.combout(\butterfly_st2[1][1][1]~1_combout ),
	.cout(\butterfly_st2[1][1][1]~2 ));
defparam \butterfly_st2[1][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][2]~1 (
	.dataa(\butterfly_st1[2][1][2]~q ),
	.datab(\butterfly_st1[3][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][1]~2 ),
	.combout(\butterfly_st2[1][1][2]~1_combout ),
	.cout(\butterfly_st2[1][1][2]~2 ));
defparam \butterfly_st2[1][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][2]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][1][10] (
	.clk(clk),
	.d(\butterfly_st1[2][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][10] .power_up = "low";

dffeas \butterfly_st1[3][0][10] (
	.clk(clk),
	.d(\butterfly_st1[3][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][10] .power_up = "low";

dffeas \butterfly_st1[2][1][9] (
	.clk(clk),
	.d(\butterfly_st1[2][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][9] .power_up = "low";

dffeas \butterfly_st1[3][0][9] (
	.clk(clk),
	.d(\butterfly_st1[3][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][9] .power_up = "low";

dffeas \butterfly_st1[2][1][8] (
	.clk(clk),
	.d(\butterfly_st1[2][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][8] .power_up = "low";

dffeas \butterfly_st1[3][0][8] (
	.clk(clk),
	.d(\butterfly_st1[3][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][8] .power_up = "low";

dffeas \butterfly_st1[2][1][7] (
	.clk(clk),
	.d(\butterfly_st1[2][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][7] .power_up = "low";

dffeas \butterfly_st1[3][0][7] (
	.clk(clk),
	.d(\butterfly_st1[3][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][7] .power_up = "low";

dffeas \butterfly_st1[2][1][6] (
	.clk(clk),
	.d(\butterfly_st1[2][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][6] .power_up = "low";

dffeas \butterfly_st1[3][0][6] (
	.clk(clk),
	.d(\butterfly_st1[3][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][6] .power_up = "low";

dffeas \butterfly_st1[2][1][5] (
	.clk(clk),
	.d(\butterfly_st1[2][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][5] .power_up = "low";

dffeas \butterfly_st1[3][0][5] (
	.clk(clk),
	.d(\butterfly_st1[3][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][5] .power_up = "low";

dffeas \butterfly_st1[2][1][4] (
	.clk(clk),
	.d(\butterfly_st1[2][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][4] .power_up = "low";

dffeas \butterfly_st1[3][0][4] (
	.clk(clk),
	.d(\butterfly_st1[3][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][4] .power_up = "low";

dffeas \butterfly_st1[2][1][3] (
	.clk(clk),
	.d(\butterfly_st1[2][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][3] .power_up = "low";

dffeas \butterfly_st1[3][0][3] (
	.clk(clk),
	.d(\butterfly_st1[3][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][3] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[1][1][3]~1 (
	.dataa(\butterfly_st1[2][1][3]~q ),
	.datab(\butterfly_st1[3][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][2]~2 ),
	.combout(\butterfly_st2[1][1][3]~1_combout ),
	.cout(\butterfly_st2[1][1][3]~2 ));
defparam \butterfly_st2[1][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][4]~1 (
	.dataa(\butterfly_st1[2][1][4]~q ),
	.datab(\butterfly_st1[3][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][3]~2 ),
	.combout(\butterfly_st2[1][1][4]~1_combout ),
	.cout(\butterfly_st2[1][1][4]~2 ));
defparam \butterfly_st2[1][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][5]~1 (
	.dataa(\butterfly_st1[2][1][5]~q ),
	.datab(\butterfly_st1[3][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][4]~2 ),
	.combout(\butterfly_st2[1][1][5]~1_combout ),
	.cout(\butterfly_st2[1][1][5]~2 ));
defparam \butterfly_st2[1][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][6]~1 (
	.dataa(\butterfly_st1[2][1][6]~q ),
	.datab(\butterfly_st1[3][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][5]~2 ),
	.combout(\butterfly_st2[1][1][6]~1_combout ),
	.cout(\butterfly_st2[1][1][6]~2 ));
defparam \butterfly_st2[1][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][7]~1 (
	.dataa(\butterfly_st1[2][1][7]~q ),
	.datab(\butterfly_st1[3][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][6]~2 ),
	.combout(\butterfly_st2[1][1][7]~1_combout ),
	.cout(\butterfly_st2[1][1][7]~2 ));
defparam \butterfly_st2[1][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][8]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][7]~2 ),
	.combout(\butterfly_st2[1][1][8]~1_combout ),
	.cout(\butterfly_st2[1][1][8]~2 ));
defparam \butterfly_st2[1][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][9]~1 (
	.dataa(\butterfly_st1[2][1][9]~q ),
	.datab(\butterfly_st1[3][0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][8]~2 ),
	.combout(\butterfly_st2[1][1][9]~1_combout ),
	.cout(\butterfly_st2[1][1][9]~2 ));
defparam \butterfly_st2[1][1][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[1][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][10]~1 (
	.dataa(\butterfly_st1[2][1][10]~q ),
	.datab(\butterfly_st1[3][0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][1][9]~2 ),
	.combout(\butterfly_st2[1][1][10]~1_combout ),
	.cout(\butterfly_st2[1][1][10]~2 ));
defparam \butterfly_st2[1][1][10]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[1][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][1][11]~1 (
	.dataa(\butterfly_st1[2][1][10]~q ),
	.datab(\butterfly_st1[3][0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[1][1][10]~2 ),
	.combout(\butterfly_st2[1][1][11]~1_combout ),
	.cout());
defparam \butterfly_st2[1][1][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[1][1][11]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][0][2] (
	.clk(clk),
	.d(\butterfly_st1[2][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][2] .power_up = "low";

dffeas \butterfly_st1[3][1][2] (
	.clk(clk),
	.d(\butterfly_st1[3][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][2] .power_up = "low";

dffeas \butterfly_st1[2][0][1] (
	.clk(clk),
	.d(\butterfly_st1[2][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][1] .power_up = "low";

dffeas \butterfly_st1[3][1][1] (
	.clk(clk),
	.d(\butterfly_st1[3][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][1] .power_up = "low";

dffeas \butterfly_st1[2][0][0] (
	.clk(clk),
	.d(\butterfly_st1[2][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][0] .power_up = "low";

dffeas \butterfly_st1[3][1][0] (
	.clk(clk),
	.d(\butterfly_st1[3][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][0] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[1][0][0]~1 (
	.dataa(\butterfly_st1[2][0][0]~q ),
	.datab(\butterfly_st1[3][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[1][0][0]~1_combout ),
	.cout(\butterfly_st2[1][0][0]~2 ));
defparam \butterfly_st2[1][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[1][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[1][0][1]~1 (
	.dataa(\butterfly_st1[2][0][1]~q ),
	.datab(\butterfly_st1[3][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][0]~2 ),
	.combout(\butterfly_st2[1][0][1]~1_combout ),
	.cout(\butterfly_st2[1][0][1]~2 ));
defparam \butterfly_st2[1][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][2]~1 (
	.dataa(\butterfly_st1[2][0][2]~q ),
	.datab(\butterfly_st1[3][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][1]~2 ),
	.combout(\butterfly_st2[1][0][2]~1_combout ),
	.cout(\butterfly_st2[1][0][2]~2 ));
defparam \butterfly_st2[1][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][2]~1 .sum_lutc_input = "cin";

dffeas \butterfly_st1[2][0][10] (
	.clk(clk),
	.d(\butterfly_st1[2][0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][10] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][10] .power_up = "low";

dffeas \butterfly_st1[3][1][10] (
	.clk(clk),
	.d(\butterfly_st1[3][1][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][10]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][10] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][10] .power_up = "low";

dffeas \butterfly_st1[2][0][9] (
	.clk(clk),
	.d(\butterfly_st1[2][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][9] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][9] .power_up = "low";

dffeas \butterfly_st1[3][1][9] (
	.clk(clk),
	.d(\butterfly_st1[3][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][9] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][9] .power_up = "low";

dffeas \butterfly_st1[2][0][8] (
	.clk(clk),
	.d(\butterfly_st1[2][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][8] .power_up = "low";

dffeas \butterfly_st1[3][1][8] (
	.clk(clk),
	.d(\butterfly_st1[3][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][8] .power_up = "low";

dffeas \butterfly_st1[2][0][7] (
	.clk(clk),
	.d(\butterfly_st1[2][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][7] .power_up = "low";

dffeas \butterfly_st1[3][1][7] (
	.clk(clk),
	.d(\butterfly_st1[3][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][7] .power_up = "low";

dffeas \butterfly_st1[2][0][6] (
	.clk(clk),
	.d(\butterfly_st1[2][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][6] .power_up = "low";

dffeas \butterfly_st1[3][1][6] (
	.clk(clk),
	.d(\butterfly_st1[3][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][6] .power_up = "low";

dffeas \butterfly_st1[2][0][5] (
	.clk(clk),
	.d(\butterfly_st1[2][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][5] .power_up = "low";

dffeas \butterfly_st1[3][1][5] (
	.clk(clk),
	.d(\butterfly_st1[3][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][5] .power_up = "low";

dffeas \butterfly_st1[2][0][4] (
	.clk(clk),
	.d(\butterfly_st1[2][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][4] .power_up = "low";

dffeas \butterfly_st1[3][1][4] (
	.clk(clk),
	.d(\butterfly_st1[3][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][4] .power_up = "low";

dffeas \butterfly_st1[2][0][3] (
	.clk(clk),
	.d(\butterfly_st1[2][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][3] .power_up = "low";

dffeas \butterfly_st1[3][1][3] (
	.clk(clk),
	.d(\butterfly_st1[3][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\butterfly_st1[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][3] .power_up = "low";

cycloneive_lcell_comb \butterfly_st2[1][0][3]~1 (
	.dataa(\butterfly_st1[2][0][3]~q ),
	.datab(\butterfly_st1[3][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][2]~2 ),
	.combout(\butterfly_st2[1][0][3]~1_combout ),
	.cout(\butterfly_st2[1][0][3]~2 ));
defparam \butterfly_st2[1][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][4]~1 (
	.dataa(\butterfly_st1[2][0][4]~q ),
	.datab(\butterfly_st1[3][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][3]~2 ),
	.combout(\butterfly_st2[1][0][4]~1_combout ),
	.cout(\butterfly_st2[1][0][4]~2 ));
defparam \butterfly_st2[1][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][5]~1 (
	.dataa(\butterfly_st1[2][0][5]~q ),
	.datab(\butterfly_st1[3][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][4]~2 ),
	.combout(\butterfly_st2[1][0][5]~1_combout ),
	.cout(\butterfly_st2[1][0][5]~2 ));
defparam \butterfly_st2[1][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][6]~1 (
	.dataa(\butterfly_st1[2][0][6]~q ),
	.datab(\butterfly_st1[3][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][5]~2 ),
	.combout(\butterfly_st2[1][0][6]~1_combout ),
	.cout(\butterfly_st2[1][0][6]~2 ));
defparam \butterfly_st2[1][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][7]~1 (
	.dataa(\butterfly_st1[2][0][7]~q ),
	.datab(\butterfly_st1[3][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][6]~2 ),
	.combout(\butterfly_st2[1][0][7]~1_combout ),
	.cout(\butterfly_st2[1][0][7]~2 ));
defparam \butterfly_st2[1][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][8]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][7]~2 ),
	.combout(\butterfly_st2[1][0][8]~1_combout ),
	.cout(\butterfly_st2[1][0][8]~2 ));
defparam \butterfly_st2[1][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][9]~1 (
	.dataa(\butterfly_st1[2][0][9]~q ),
	.datab(\butterfly_st1[3][1][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][8]~2 ),
	.combout(\butterfly_st2[1][0][9]~1_combout ),
	.cout(\butterfly_st2[1][0][9]~2 ));
defparam \butterfly_st2[1][0][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[1][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][10]~1 (
	.dataa(\butterfly_st1[2][0][10]~q ),
	.datab(\butterfly_st1[3][1][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[1][0][9]~2 ),
	.combout(\butterfly_st2[1][0][10]~1_combout ),
	.cout(\butterfly_st2[1][0][10]~2 ));
defparam \butterfly_st2[1][0][10]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[1][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[1][0][11]~1 (
	.dataa(\butterfly_st1[2][0][10]~q ),
	.datab(\butterfly_st1[3][1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[1][0][10]~2 ),
	.combout(\butterfly_st2[1][0][11]~1_combout ),
	.cout());
defparam \butterfly_st2[1][0][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[1][0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][0]~1 (
	.dataa(\butterfly_st1[0][1][0]~q ),
	.datab(\butterfly_st1[1][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[2][1][0]~1_combout ),
	.cout(\butterfly_st2[2][1][0]~2 ));
defparam \butterfly_st2[2][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[2][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[2][1][1]~1 (
	.dataa(\butterfly_st1[0][1][1]~q ),
	.datab(\butterfly_st1[1][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][0]~2 ),
	.combout(\butterfly_st2[2][1][1]~1_combout ),
	.cout(\butterfly_st2[2][1][1]~2 ));
defparam \butterfly_st2[2][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][2]~1 (
	.dataa(\butterfly_st1[0][1][2]~q ),
	.datab(\butterfly_st1[1][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][1]~2 ),
	.combout(\butterfly_st2[2][1][2]~1_combout ),
	.cout(\butterfly_st2[2][1][2]~2 ));
defparam \butterfly_st2[2][1][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][3]~1 (
	.dataa(\butterfly_st1[0][1][3]~q ),
	.datab(\butterfly_st1[1][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][2]~2 ),
	.combout(\butterfly_st2[2][1][3]~1_combout ),
	.cout(\butterfly_st2[2][1][3]~2 ));
defparam \butterfly_st2[2][1][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][4]~1 (
	.dataa(\butterfly_st1[0][1][4]~q ),
	.datab(\butterfly_st1[1][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][3]~2 ),
	.combout(\butterfly_st2[2][1][4]~1_combout ),
	.cout(\butterfly_st2[2][1][4]~2 ));
defparam \butterfly_st2[2][1][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][5]~1 (
	.dataa(\butterfly_st1[0][1][5]~q ),
	.datab(\butterfly_st1[1][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][4]~2 ),
	.combout(\butterfly_st2[2][1][5]~1_combout ),
	.cout(\butterfly_st2[2][1][5]~2 ));
defparam \butterfly_st2[2][1][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][6]~1 (
	.dataa(\butterfly_st1[0][1][6]~q ),
	.datab(\butterfly_st1[1][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][5]~2 ),
	.combout(\butterfly_st2[2][1][6]~1_combout ),
	.cout(\butterfly_st2[2][1][6]~2 ));
defparam \butterfly_st2[2][1][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][7]~1 (
	.dataa(\butterfly_st1[0][1][7]~q ),
	.datab(\butterfly_st1[1][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][6]~2 ),
	.combout(\butterfly_st2[2][1][7]~1_combout ),
	.cout(\butterfly_st2[2][1][7]~2 ));
defparam \butterfly_st2[2][1][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][8]~1 (
	.dataa(\butterfly_st1[0][1][8]~q ),
	.datab(\butterfly_st1[1][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][7]~2 ),
	.combout(\butterfly_st2[2][1][8]~1_combout ),
	.cout(\butterfly_st2[2][1][8]~2 ));
defparam \butterfly_st2[2][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][9]~1 (
	.dataa(\butterfly_st1[0][1][9]~q ),
	.datab(\butterfly_st1[1][1][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][8]~2 ),
	.combout(\butterfly_st2[2][1][9]~1_combout ),
	.cout(\butterfly_st2[2][1][9]~2 ));
defparam \butterfly_st2[2][1][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][10]~1 (
	.dataa(\butterfly_st1[0][1][10]~q ),
	.datab(\butterfly_st1[1][1][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][1][9]~2 ),
	.combout(\butterfly_st2[2][1][10]~1_combout ),
	.cout(\butterfly_st2[2][1][10]~2 ));
defparam \butterfly_st2[2][1][10]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][1][11]~1 (
	.dataa(\butterfly_st1[0][1][10]~q ),
	.datab(\butterfly_st1[1][1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[2][1][10]~2 ),
	.combout(\butterfly_st2[2][1][11]~1_combout ),
	.cout());
defparam \butterfly_st2[2][1][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[2][1][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][0]~1 (
	.dataa(\butterfly_st1[0][0][0]~q ),
	.datab(\butterfly_st1[1][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[2][0][0]~1_combout ),
	.cout(\butterfly_st2[2][0][0]~2 ));
defparam \butterfly_st2[2][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[2][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[2][0][1]~1 (
	.dataa(\butterfly_st1[0][0][1]~q ),
	.datab(\butterfly_st1[1][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][0]~2 ),
	.combout(\butterfly_st2[2][0][1]~1_combout ),
	.cout(\butterfly_st2[2][0][1]~2 ));
defparam \butterfly_st2[2][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][2]~1 (
	.dataa(\butterfly_st1[0][0][2]~q ),
	.datab(\butterfly_st1[1][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][1]~2 ),
	.combout(\butterfly_st2[2][0][2]~1_combout ),
	.cout(\butterfly_st2[2][0][2]~2 ));
defparam \butterfly_st2[2][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][3]~1 (
	.dataa(\butterfly_st1[0][0][3]~q ),
	.datab(\butterfly_st1[1][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][2]~2 ),
	.combout(\butterfly_st2[2][0][3]~1_combout ),
	.cout(\butterfly_st2[2][0][3]~2 ));
defparam \butterfly_st2[2][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][4]~1 (
	.dataa(\butterfly_st1[0][0][4]~q ),
	.datab(\butterfly_st1[1][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][3]~2 ),
	.combout(\butterfly_st2[2][0][4]~1_combout ),
	.cout(\butterfly_st2[2][0][4]~2 ));
defparam \butterfly_st2[2][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][5]~1 (
	.dataa(\butterfly_st1[0][0][5]~q ),
	.datab(\butterfly_st1[1][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][4]~2 ),
	.combout(\butterfly_st2[2][0][5]~1_combout ),
	.cout(\butterfly_st2[2][0][5]~2 ));
defparam \butterfly_st2[2][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][6]~1 (
	.dataa(\butterfly_st1[0][0][6]~q ),
	.datab(\butterfly_st1[1][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][5]~2 ),
	.combout(\butterfly_st2[2][0][6]~1_combout ),
	.cout(\butterfly_st2[2][0][6]~2 ));
defparam \butterfly_st2[2][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][7]~1 (
	.dataa(\butterfly_st1[0][0][7]~q ),
	.datab(\butterfly_st1[1][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][6]~2 ),
	.combout(\butterfly_st2[2][0][7]~1_combout ),
	.cout(\butterfly_st2[2][0][7]~2 ));
defparam \butterfly_st2[2][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][8]~1 (
	.dataa(\butterfly_st1[0][0][8]~q ),
	.datab(\butterfly_st1[1][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][7]~2 ),
	.combout(\butterfly_st2[2][0][8]~1_combout ),
	.cout(\butterfly_st2[2][0][8]~2 ));
defparam \butterfly_st2[2][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][9]~1 (
	.dataa(\butterfly_st1[0][0][9]~q ),
	.datab(\butterfly_st1[1][0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][8]~2 ),
	.combout(\butterfly_st2[2][0][9]~1_combout ),
	.cout(\butterfly_st2[2][0][9]~2 ));
defparam \butterfly_st2[2][0][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[2][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][10]~1 (
	.dataa(\butterfly_st1[0][0][10]~q ),
	.datab(\butterfly_st1[1][0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[2][0][9]~2 ),
	.combout(\butterfly_st2[2][0][10]~1_combout ),
	.cout(\butterfly_st2[2][0][10]~2 ));
defparam \butterfly_st2[2][0][10]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[2][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[2][0][11]~1 (
	.dataa(\butterfly_st1[0][0][10]~q ),
	.datab(\butterfly_st1[1][0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[2][0][10]~2 ),
	.combout(\butterfly_st2[2][0][11]~1_combout ),
	.cout());
defparam \butterfly_st2[2][0][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[2][0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][0]~1 (
	.dataa(\butterfly_st1[2][1][0]~q ),
	.datab(\butterfly_st1[3][0][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[3][1][0]~1_combout ),
	.cout(\butterfly_st2[3][1][0]~2 ));
defparam \butterfly_st2[3][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st2[3][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[3][1][1]~1 (
	.dataa(\butterfly_st1[2][1][1]~q ),
	.datab(\butterfly_st1[3][0][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][0]~2 ),
	.combout(\butterfly_st2[3][1][1]~1_combout ),
	.cout(\butterfly_st2[3][1][1]~2 ));
defparam \butterfly_st2[3][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][2]~1 (
	.dataa(\butterfly_st1[2][1][2]~q ),
	.datab(\butterfly_st1[3][0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][1]~2 ),
	.combout(\butterfly_st2[3][1][2]~1_combout ),
	.cout(\butterfly_st2[3][1][2]~2 ));
defparam \butterfly_st2[3][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][3]~1 (
	.dataa(\butterfly_st1[2][1][3]~q ),
	.datab(\butterfly_st1[3][0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][2]~2 ),
	.combout(\butterfly_st2[3][1][3]~1_combout ),
	.cout(\butterfly_st2[3][1][3]~2 ));
defparam \butterfly_st2[3][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][4]~1 (
	.dataa(\butterfly_st1[2][1][4]~q ),
	.datab(\butterfly_st1[3][0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][3]~2 ),
	.combout(\butterfly_st2[3][1][4]~1_combout ),
	.cout(\butterfly_st2[3][1][4]~2 ));
defparam \butterfly_st2[3][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][5]~1 (
	.dataa(\butterfly_st1[2][1][5]~q ),
	.datab(\butterfly_st1[3][0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][4]~2 ),
	.combout(\butterfly_st2[3][1][5]~1_combout ),
	.cout(\butterfly_st2[3][1][5]~2 ));
defparam \butterfly_st2[3][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][6]~1 (
	.dataa(\butterfly_st1[2][1][6]~q ),
	.datab(\butterfly_st1[3][0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][5]~2 ),
	.combout(\butterfly_st2[3][1][6]~1_combout ),
	.cout(\butterfly_st2[3][1][6]~2 ));
defparam \butterfly_st2[3][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][7]~1 (
	.dataa(\butterfly_st1[2][1][7]~q ),
	.datab(\butterfly_st1[3][0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][6]~2 ),
	.combout(\butterfly_st2[3][1][7]~1_combout ),
	.cout(\butterfly_st2[3][1][7]~2 ));
defparam \butterfly_st2[3][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][8]~1 (
	.dataa(\butterfly_st1[2][1][8]~q ),
	.datab(\butterfly_st1[3][0][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][7]~2 ),
	.combout(\butterfly_st2[3][1][8]~1_combout ),
	.cout(\butterfly_st2[3][1][8]~2 ));
defparam \butterfly_st2[3][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][9]~1 (
	.dataa(\butterfly_st1[2][1][9]~q ),
	.datab(\butterfly_st1[3][0][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][8]~2 ),
	.combout(\butterfly_st2[3][1][9]~1_combout ),
	.cout(\butterfly_st2[3][1][9]~2 ));
defparam \butterfly_st2[3][1][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st2[3][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][10]~1 (
	.dataa(\butterfly_st1[2][1][10]~q ),
	.datab(\butterfly_st1[3][0][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][1][9]~2 ),
	.combout(\butterfly_st2[3][1][10]~1_combout ),
	.cout(\butterfly_st2[3][1][10]~2 ));
defparam \butterfly_st2[3][1][10]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st2[3][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][1][11]~1 (
	.dataa(\butterfly_st1[2][1][10]~q ),
	.datab(\butterfly_st1[3][0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[3][1][10]~2 ),
	.combout(\butterfly_st2[3][1][11]~1_combout ),
	.cout());
defparam \butterfly_st2[3][1][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[3][1][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][0]~1 (
	.dataa(\butterfly_st1[2][0][0]~q ),
	.datab(\butterfly_st1[3][1][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st2[3][0][0]~1_combout ),
	.cout(\butterfly_st2[3][0][0]~2 ));
defparam \butterfly_st2[3][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st2[3][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st2[3][0][1]~1 (
	.dataa(\butterfly_st1[2][0][1]~q ),
	.datab(\butterfly_st1[3][1][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][0]~2 ),
	.combout(\butterfly_st2[3][0][1]~1_combout ),
	.cout(\butterfly_st2[3][0][1]~2 ));
defparam \butterfly_st2[3][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][2]~1 (
	.dataa(\butterfly_st1[2][0][2]~q ),
	.datab(\butterfly_st1[3][1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][1]~2 ),
	.combout(\butterfly_st2[3][0][2]~1_combout ),
	.cout(\butterfly_st2[3][0][2]~2 ));
defparam \butterfly_st2[3][0][2]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][3]~1 (
	.dataa(\butterfly_st1[2][0][3]~q ),
	.datab(\butterfly_st1[3][1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][2]~2 ),
	.combout(\butterfly_st2[3][0][3]~1_combout ),
	.cout(\butterfly_st2[3][0][3]~2 ));
defparam \butterfly_st2[3][0][3]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][4]~1 (
	.dataa(\butterfly_st1[2][0][4]~q ),
	.datab(\butterfly_st1[3][1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][3]~2 ),
	.combout(\butterfly_st2[3][0][4]~1_combout ),
	.cout(\butterfly_st2[3][0][4]~2 ));
defparam \butterfly_st2[3][0][4]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][5]~1 (
	.dataa(\butterfly_st1[2][0][5]~q ),
	.datab(\butterfly_st1[3][1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][4]~2 ),
	.combout(\butterfly_st2[3][0][5]~1_combout ),
	.cout(\butterfly_st2[3][0][5]~2 ));
defparam \butterfly_st2[3][0][5]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][6]~1 (
	.dataa(\butterfly_st1[2][0][6]~q ),
	.datab(\butterfly_st1[3][1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][5]~2 ),
	.combout(\butterfly_st2[3][0][6]~1_combout ),
	.cout(\butterfly_st2[3][0][6]~2 ));
defparam \butterfly_st2[3][0][6]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][7]~1 (
	.dataa(\butterfly_st1[2][0][7]~q ),
	.datab(\butterfly_st1[3][1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][6]~2 ),
	.combout(\butterfly_st2[3][0][7]~1_combout ),
	.cout(\butterfly_st2[3][0][7]~2 ));
defparam \butterfly_st2[3][0][7]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][8]~1 (
	.dataa(\butterfly_st1[2][0][8]~q ),
	.datab(\butterfly_st1[3][1][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][7]~2 ),
	.combout(\butterfly_st2[3][0][8]~1_combout ),
	.cout(\butterfly_st2[3][0][8]~2 ));
defparam \butterfly_st2[3][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][9]~1 (
	.dataa(\butterfly_st1[2][0][9]~q ),
	.datab(\butterfly_st1[3][1][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][8]~2 ),
	.combout(\butterfly_st2[3][0][9]~1_combout ),
	.cout(\butterfly_st2[3][0][9]~2 ));
defparam \butterfly_st2[3][0][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st2[3][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][10]~1 (
	.dataa(\butterfly_st1[2][0][10]~q ),
	.datab(\butterfly_st1[3][1][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st2[3][0][9]~2 ),
	.combout(\butterfly_st2[3][0][10]~1_combout ),
	.cout(\butterfly_st2[3][0][10]~2 ));
defparam \butterfly_st2[3][0][10]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st2[3][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st2[3][0][11]~1 (
	.dataa(\butterfly_st1[2][0][10]~q ),
	.datab(\butterfly_st1[3][1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st2[3][0][10]~2 ),
	.combout(\butterfly_st2[3][0][11]~1_combout ),
	.cout());
defparam \butterfly_st2[3][0][11]~1 .lut_mask = 16'h9696;
defparam \butterfly_st2[3][0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][0]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[0][0][0]~1_combout ),
	.cout(\butterfly_st1[0][0][0]~2 ));
defparam \butterfly_st1[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[0][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[0][0][1]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][0]~2 ),
	.combout(\butterfly_st1[0][0][1]~1_combout ),
	.cout(\butterfly_st1[0][0][1]~2 ));
defparam \butterfly_st1[0][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][2]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][1]~2 ),
	.combout(\butterfly_st1[0][0][2]~1_combout ),
	.cout(\butterfly_st1[0][0][2]~2 ));
defparam \butterfly_st1[0][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][3]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][2]~2 ),
	.combout(\butterfly_st1[0][0][3]~1_combout ),
	.cout(\butterfly_st1[0][0][3]~2 ));
defparam \butterfly_st1[0][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][4]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][3]~2 ),
	.combout(\butterfly_st1[0][0][4]~1_combout ),
	.cout(\butterfly_st1[0][0][4]~2 ));
defparam \butterfly_st1[0][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][5]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][4]~2 ),
	.combout(\butterfly_st1[0][0][5]~1_combout ),
	.cout(\butterfly_st1[0][0][5]~2 ));
defparam \butterfly_st1[0][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][6]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][5]~2 ),
	.combout(\butterfly_st1[0][0][6]~1_combout ),
	.cout(\butterfly_st1[0][0][6]~2 ));
defparam \butterfly_st1[0][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][7]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][6]~2 ),
	.combout(\butterfly_st1[0][0][7]~1_combout ),
	.cout(\butterfly_st1[0][0][7]~2 ));
defparam \butterfly_st1[0][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][8]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][8]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][7]~2 ),
	.combout(\butterfly_st1[0][0][8]~1_combout ),
	.cout(\butterfly_st1[0][0][8]~2 ));
defparam \butterfly_st1[0][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][0]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[1][0][0]~1_combout ),
	.cout(\butterfly_st1[1][0][0]~2 ));
defparam \butterfly_st1[1][0][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[1][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[1][0][1]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][0]~2 ),
	.combout(\butterfly_st1[1][0][1]~1_combout ),
	.cout(\butterfly_st1[1][0][1]~2 ));
defparam \butterfly_st1[1][0][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][2]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][1]~2 ),
	.combout(\butterfly_st1[1][0][2]~1_combout ),
	.cout(\butterfly_st1[1][0][2]~2 ));
defparam \butterfly_st1[1][0][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][3]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][2]~2 ),
	.combout(\butterfly_st1[1][0][3]~1_combout ),
	.cout(\butterfly_st1[1][0][3]~2 ));
defparam \butterfly_st1[1][0][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][4]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][3]~2 ),
	.combout(\butterfly_st1[1][0][4]~1_combout ),
	.cout(\butterfly_st1[1][0][4]~2 ));
defparam \butterfly_st1[1][0][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][5]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][4]~2 ),
	.combout(\butterfly_st1[1][0][5]~1_combout ),
	.cout(\butterfly_st1[1][0][5]~2 ));
defparam \butterfly_st1[1][0][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][6]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][5]~2 ),
	.combout(\butterfly_st1[1][0][6]~1_combout ),
	.cout(\butterfly_st1[1][0][6]~2 ));
defparam \butterfly_st1[1][0][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][7]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][6]~2 ),
	.combout(\butterfly_st1[1][0][7]~1_combout ),
	.cout(\butterfly_st1[1][0][7]~2 ));
defparam \butterfly_st1[1][0][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][8]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][8]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][7]~2 ),
	.combout(\butterfly_st1[1][0][8]~1_combout ),
	.cout(\butterfly_st1[1][0][8]~2 ));
defparam \butterfly_st1[1][0][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][9]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][0][8]~2 ),
	.combout(\butterfly_st1[0][0][9]~1_combout ),
	.cout(\butterfly_st1[0][0][9]~2 ));
defparam \butterfly_st1[0][0][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][0][10]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[0][0][9]~2 ),
	.combout(\butterfly_st1[0][0][10]~1_combout ),
	.cout());
defparam \butterfly_st1[0][0][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[0][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][9]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][0][8]~2 ),
	.combout(\butterfly_st1[1][0][9]~1_combout ),
	.cout(\butterfly_st1[1][0][9]~2 ));
defparam \butterfly_st1[1][0][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][0][10]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[1][0][9]~2 ),
	.combout(\butterfly_st1[1][0][10]~1_combout ),
	.cout());
defparam \butterfly_st1[1][0][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[1][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][0]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[0][1][0]~1_combout ),
	.cout(\butterfly_st1[0][1][0]~2 ));
defparam \butterfly_st1[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[0][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[0][1][1]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][0]~2 ),
	.combout(\butterfly_st1[0][1][1]~1_combout ),
	.cout(\butterfly_st1[0][1][1]~2 ));
defparam \butterfly_st1[0][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][2]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][1]~2 ),
	.combout(\butterfly_st1[0][1][2]~1_combout ),
	.cout(\butterfly_st1[0][1][2]~2 ));
defparam \butterfly_st1[0][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][3]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][2]~2 ),
	.combout(\butterfly_st1[0][1][3]~1_combout ),
	.cout(\butterfly_st1[0][1][3]~2 ));
defparam \butterfly_st1[0][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][4]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][3]~2 ),
	.combout(\butterfly_st1[0][1][4]~1_combout ),
	.cout(\butterfly_st1[0][1][4]~2 ));
defparam \butterfly_st1[0][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][5]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][4]~2 ),
	.combout(\butterfly_st1[0][1][5]~1_combout ),
	.cout(\butterfly_st1[0][1][5]~2 ));
defparam \butterfly_st1[0][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][6]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][5]~2 ),
	.combout(\butterfly_st1[0][1][6]~1_combout ),
	.cout(\butterfly_st1[0][1][6]~2 ));
defparam \butterfly_st1[0][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][7]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][6]~2 ),
	.combout(\butterfly_st1[0][1][7]~1_combout ),
	.cout(\butterfly_st1[0][1][7]~2 ));
defparam \butterfly_st1[0][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][8]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][8]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][7]~2 ),
	.combout(\butterfly_st1[0][1][8]~1_combout ),
	.cout(\butterfly_st1[0][1][8]~2 ));
defparam \butterfly_st1[0][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[0][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][0]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[1][1][0]~1_combout ),
	.cout(\butterfly_st1[1][1][0]~2 ));
defparam \butterfly_st1[1][1][0]~1 .lut_mask = 16'h66EE;
defparam \butterfly_st1[1][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[1][1][1]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][0]~2 ),
	.combout(\butterfly_st1[1][1][1]~1_combout ),
	.cout(\butterfly_st1[1][1][1]~2 ));
defparam \butterfly_st1[1][1][1]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][2]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][1]~2 ),
	.combout(\butterfly_st1[1][1][2]~1_combout ),
	.cout(\butterfly_st1[1][1][2]~2 ));
defparam \butterfly_st1[1][1][2]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][3]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][2]~2 ),
	.combout(\butterfly_st1[1][1][3]~1_combout ),
	.cout(\butterfly_st1[1][1][3]~2 ));
defparam \butterfly_st1[1][1][3]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][4]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][3]~2 ),
	.combout(\butterfly_st1[1][1][4]~1_combout ),
	.cout(\butterfly_st1[1][1][4]~2 ));
defparam \butterfly_st1[1][1][4]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][5]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][4]~2 ),
	.combout(\butterfly_st1[1][1][5]~1_combout ),
	.cout(\butterfly_st1[1][1][5]~2 ));
defparam \butterfly_st1[1][1][5]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][6]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][5]~2 ),
	.combout(\butterfly_st1[1][1][6]~1_combout ),
	.cout(\butterfly_st1[1][1][6]~2 ));
defparam \butterfly_st1[1][1][6]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][7]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][6]~2 ),
	.combout(\butterfly_st1[1][1][7]~1_combout ),
	.cout(\butterfly_st1[1][1][7]~2 ));
defparam \butterfly_st1[1][1][7]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][8]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][8]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][7]~2 ),
	.combout(\butterfly_st1[1][1][8]~1_combout ),
	.cout(\butterfly_st1[1][1][8]~2 ));
defparam \butterfly_st1[1][1][8]~1 .lut_mask = 16'h96EF;
defparam \butterfly_st1[1][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][9]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[0][1][8]~2 ),
	.combout(\butterfly_st1[0][1][9]~1_combout ),
	.cout(\butterfly_st1[0][1][9]~2 ));
defparam \butterfly_st1[0][1][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[0][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[0][1][10]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[0][1][9]~2 ),
	.combout(\butterfly_st1[0][1][10]~1_combout ),
	.cout());
defparam \butterfly_st1[0][1][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[0][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][9]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[1][1][8]~2 ),
	.combout(\butterfly_st1[1][1][9]~1_combout ),
	.cout(\butterfly_st1[1][1][9]~2 ));
defparam \butterfly_st1[1][1][9]~1 .lut_mask = 16'h967F;
defparam \butterfly_st1[1][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[1][1][10]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[1][1][9]~2 ),
	.combout(\butterfly_st1[1][1][10]~1_combout ),
	.cout());
defparam \butterfly_st1[1][1][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[1][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][0]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[2][1][0]~1_combout ),
	.cout(\butterfly_st1[2][1][0]~2 ));
defparam \butterfly_st1[2][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[2][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[2][1][1]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][0]~2 ),
	.combout(\butterfly_st1[2][1][1]~1_combout ),
	.cout(\butterfly_st1[2][1][1]~2 ));
defparam \butterfly_st1[2][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][2]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][1]~2 ),
	.combout(\butterfly_st1[2][1][2]~1_combout ),
	.cout(\butterfly_st1[2][1][2]~2 ));
defparam \butterfly_st1[2][1][2]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][0]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[3][0][0]~1_combout ),
	.cout(\butterfly_st1[3][0][0]~2 ));
defparam \butterfly_st1[3][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[3][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[3][0][1]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][0]~2 ),
	.combout(\butterfly_st1[3][0][1]~1_combout ),
	.cout(\butterfly_st1[3][0][1]~2 ));
defparam \butterfly_st1[3][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][2]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][1]~2 ),
	.combout(\butterfly_st1[3][0][2]~1_combout ),
	.cout(\butterfly_st1[3][0][2]~2 ));
defparam \butterfly_st1[3][0][2]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][3]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][2]~2 ),
	.combout(\butterfly_st1[2][1][3]~1_combout ),
	.cout(\butterfly_st1[2][1][3]~2 ));
defparam \butterfly_st1[2][1][3]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][4]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][3]~2 ),
	.combout(\butterfly_st1[2][1][4]~1_combout ),
	.cout(\butterfly_st1[2][1][4]~2 ));
defparam \butterfly_st1[2][1][4]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][5]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][4]~2 ),
	.combout(\butterfly_st1[2][1][5]~1_combout ),
	.cout(\butterfly_st1[2][1][5]~2 ));
defparam \butterfly_st1[2][1][5]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][6]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][5]~2 ),
	.combout(\butterfly_st1[2][1][6]~1_combout ),
	.cout(\butterfly_st1[2][1][6]~2 ));
defparam \butterfly_st1[2][1][6]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][7]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][6]~2 ),
	.combout(\butterfly_st1[2][1][7]~1_combout ),
	.cout(\butterfly_st1[2][1][7]~2 ));
defparam \butterfly_st1[2][1][7]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][8]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][8]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][7]~2 ),
	.combout(\butterfly_st1[2][1][8]~1_combout ),
	.cout(\butterfly_st1[2][1][8]~2 ));
defparam \butterfly_st1[2][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][9]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][1][8]~2 ),
	.combout(\butterfly_st1[2][1][9]~1_combout ),
	.cout(\butterfly_st1[2][1][9]~2 ));
defparam \butterfly_st1[2][1][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][1][10]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[2][1][9]~2 ),
	.combout(\butterfly_st1[2][1][10]~1_combout ),
	.cout());
defparam \butterfly_st1[2][1][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[2][1][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][3]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][2]~2 ),
	.combout(\butterfly_st1[3][0][3]~1_combout ),
	.cout(\butterfly_st1[3][0][3]~2 ));
defparam \butterfly_st1[3][0][3]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][4]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][3]~2 ),
	.combout(\butterfly_st1[3][0][4]~1_combout ),
	.cout(\butterfly_st1[3][0][4]~2 ));
defparam \butterfly_st1[3][0][4]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][5]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][4]~2 ),
	.combout(\butterfly_st1[3][0][5]~1_combout ),
	.cout(\butterfly_st1[3][0][5]~2 ));
defparam \butterfly_st1[3][0][5]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][6]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][5]~2 ),
	.combout(\butterfly_st1[3][0][6]~1_combout ),
	.cout(\butterfly_st1[3][0][6]~2 ));
defparam \butterfly_st1[3][0][6]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][7]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][6]~2 ),
	.combout(\butterfly_st1[3][0][7]~1_combout ),
	.cout(\butterfly_st1[3][0][7]~2 ));
defparam \butterfly_st1[3][0][7]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][8]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][8]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][7]~2 ),
	.combout(\butterfly_st1[3][0][8]~1_combout ),
	.cout(\butterfly_st1[3][0][8]~2 ));
defparam \butterfly_st1[3][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][9]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][0][8]~2 ),
	.combout(\butterfly_st1[3][0][9]~1_combout ),
	.cout(\butterfly_st1[3][0][9]~2 ));
defparam \butterfly_st1[3][0][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][0][10]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[3][0][9]~2 ),
	.combout(\butterfly_st1[3][0][10]~1_combout ),
	.cout());
defparam \butterfly_st1[3][0][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[3][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][0]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[2][0][0]~1_combout ),
	.cout(\butterfly_st1[2][0][0]~2 ));
defparam \butterfly_st1[2][0][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[2][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[2][0][1]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][0]~2 ),
	.combout(\butterfly_st1[2][0][1]~1_combout ),
	.cout(\butterfly_st1[2][0][1]~2 ));
defparam \butterfly_st1[2][0][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][2]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][1]~2 ),
	.combout(\butterfly_st1[2][0][2]~1_combout ),
	.cout(\butterfly_st1[2][0][2]~2 ));
defparam \butterfly_st1[2][0][2]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][0]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\butterfly_st1[3][1][0]~1_combout ),
	.cout(\butterfly_st1[3][1][0]~2 ));
defparam \butterfly_st1[3][1][0]~1 .lut_mask = 16'h66BB;
defparam \butterfly_st1[3][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \butterfly_st1[3][1][1]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][0]~2 ),
	.combout(\butterfly_st1[3][1][1]~1_combout ),
	.cout(\butterfly_st1[3][1][1]~2 ));
defparam \butterfly_st1[3][1][1]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][2]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][1]~2 ),
	.combout(\butterfly_st1[3][1][2]~1_combout ),
	.cout(\butterfly_st1[3][1][2]~2 ));
defparam \butterfly_st1[3][1][2]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][3]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][2]~2 ),
	.combout(\butterfly_st1[2][0][3]~1_combout ),
	.cout(\butterfly_st1[2][0][3]~2 ));
defparam \butterfly_st1[2][0][3]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][4]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][3]~2 ),
	.combout(\butterfly_st1[2][0][4]~1_combout ),
	.cout(\butterfly_st1[2][0][4]~2 ));
defparam \butterfly_st1[2][0][4]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][5]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][4]~2 ),
	.combout(\butterfly_st1[2][0][5]~1_combout ),
	.cout(\butterfly_st1[2][0][5]~2 ));
defparam \butterfly_st1[2][0][5]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][6]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][5]~2 ),
	.combout(\butterfly_st1[2][0][6]~1_combout ),
	.cout(\butterfly_st1[2][0][6]~2 ));
defparam \butterfly_st1[2][0][6]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][7]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][6]~2 ),
	.combout(\butterfly_st1[2][0][7]~1_combout ),
	.cout(\butterfly_st1[2][0][7]~2 ));
defparam \butterfly_st1[2][0][7]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][8]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][8]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][7]~2 ),
	.combout(\butterfly_st1[2][0][8]~1_combout ),
	.cout(\butterfly_st1[2][0][8]~2 ));
defparam \butterfly_st1[2][0][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[2][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][9]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[2][0][8]~2 ),
	.combout(\butterfly_st1[2][0][9]~1_combout ),
	.cout(\butterfly_st1[2][0][9]~2 ));
defparam \butterfly_st1[2][0][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[2][0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[2][0][10]~1 (
	.dataa(\gen_disc:bfp_scale|r_array_out[0][9]~q ),
	.datab(\gen_disc:bfp_scale|r_array_out[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[2][0][9]~2 ),
	.combout(\butterfly_st1[2][0][10]~1_combout ),
	.cout());
defparam \butterfly_st1[2][0][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[2][0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][3]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][2]~2 ),
	.combout(\butterfly_st1[3][1][3]~1_combout ),
	.cout(\butterfly_st1[3][1][3]~2 ));
defparam \butterfly_st1[3][1][3]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][4]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][3]~2 ),
	.combout(\butterfly_st1[3][1][4]~1_combout ),
	.cout(\butterfly_st1[3][1][4]~2 ));
defparam \butterfly_st1[3][1][4]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][5]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][4]~2 ),
	.combout(\butterfly_st1[3][1][5]~1_combout ),
	.cout(\butterfly_st1[3][1][5]~2 ));
defparam \butterfly_st1[3][1][5]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][6]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][5]~2 ),
	.combout(\butterfly_st1[3][1][6]~1_combout ),
	.cout(\butterfly_st1[3][1][6]~2 ));
defparam \butterfly_st1[3][1][6]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][7]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][6]~2 ),
	.combout(\butterfly_st1[3][1][7]~1_combout ),
	.cout(\butterfly_st1[3][1][7]~2 ));
defparam \butterfly_st1[3][1][7]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][8]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][8]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][7]~2 ),
	.combout(\butterfly_st1[3][1][8]~1_combout ),
	.cout(\butterfly_st1[3][1][8]~2 ));
defparam \butterfly_st1[3][1][8]~1 .lut_mask = 16'h96BF;
defparam \butterfly_st1[3][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][9]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\butterfly_st1[3][1][8]~2 ),
	.combout(\butterfly_st1[3][1][9]~1_combout ),
	.cout(\butterfly_st1[3][1][9]~2 ));
defparam \butterfly_st1[3][1][9]~1 .lut_mask = 16'h96DF;
defparam \butterfly_st1[3][1][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \butterfly_st1[3][1][10]~1 (
	.dataa(\gen_disc:bfp_scale|i_array_out[1][9]~q ),
	.datab(\gen_disc:bfp_scale|i_array_out[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\butterfly_st1[3][1][9]~2 ),
	.combout(\butterfly_st1[3][1][10]~1_combout ),
	.cout());
defparam \butterfly_st1[3][1][10]~1 .lut_mask = 16'h9696;
defparam \butterfly_st1[3][1][10]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[6][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle605),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][5] .power_up = "low";

dffeas \reg_no_twiddle[6][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle609),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][9] .power_up = "low";

dffeas \reg_no_twiddle[6][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle615),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][5] .power_up = "low";

dffeas \reg_no_twiddle[6][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle619),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][9] .power_up = "low";

dffeas \reg_no_twiddle[6][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle606),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][6] .power_up = "low";

dffeas \reg_no_twiddle[6][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle616),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][6] .power_up = "low";

dffeas \reg_no_twiddle[6][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle607),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][7] .power_up = "low";

dffeas \reg_no_twiddle[6][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle617),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][7] .power_up = "low";

dffeas \reg_no_twiddle[6][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle608),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][8] .power_up = "low";

dffeas \reg_no_twiddle[6][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle618),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][8] .power_up = "low";

dffeas \reg_no_twiddle[6][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle602),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][2] .power_up = "low";

dffeas \reg_no_twiddle[6][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle612),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][2] .power_up = "low";

dffeas \reg_no_twiddle[6][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle601),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][1] .power_up = "low";

dffeas \reg_no_twiddle[6][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle611),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][1] .power_up = "low";

dffeas \reg_no_twiddle[6][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle600),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][0] .power_up = "low";

dffeas \reg_no_twiddle[6][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle610),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][0] .power_up = "low";

dffeas \reg_no_twiddle[6][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle604),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][4] .power_up = "low";

dffeas \reg_no_twiddle[6][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle614),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][4] .power_up = "low";

dffeas \reg_no_twiddle[6][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle603),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][3] .power_up = "low";

dffeas \reg_no_twiddle[6][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(reg_no_twiddle613),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~80 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.cin(gnd),
	.combout(\reg_no_twiddle~80_combout ),
	.cout());
defparam \reg_no_twiddle~80 .lut_mask = 16'hAAFF;
defparam \reg_no_twiddle~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][0][0]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\reg_no_twiddle~80_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\reg_no_twiddle[0][0][0]~1_combout ),
	.cout(\reg_no_twiddle[0][0][0]~2 ));
defparam \reg_no_twiddle[0][0][0]~1 .lut_mask = 16'h66EE;
defparam \reg_no_twiddle[0][0][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][0][1]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][0]~2 ),
	.combout(\reg_no_twiddle[0][0][1]~1_combout ),
	.cout(\reg_no_twiddle[0][0][1]~2 ));
defparam \reg_no_twiddle[0][0][1]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][2]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][1]~2 ),
	.combout(\reg_no_twiddle[0][0][2]~1_combout ),
	.cout(\reg_no_twiddle[0][0][2]~2 ));
defparam \reg_no_twiddle[0][0][2]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][3]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][2]~2 ),
	.combout(\reg_no_twiddle[0][0][3]~1_combout ),
	.cout(\reg_no_twiddle[0][0][3]~2 ));
defparam \reg_no_twiddle[0][0][3]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][4]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][3]~2 ),
	.combout(\reg_no_twiddle[0][0][4]~1_combout ),
	.cout(\reg_no_twiddle[0][0][4]~2 ));
defparam \reg_no_twiddle[0][0][4]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][5]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][4]~2 ),
	.combout(\reg_no_twiddle[0][0][5]~1_combout ),
	.cout(\reg_no_twiddle[0][0][5]~2 ));
defparam \reg_no_twiddle[0][0][5]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][5]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~60 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~60_combout ),
	.cout());
defparam \reg_no_twiddle~60 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~60 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~40 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~40_combout ),
	.cout());
defparam \reg_no_twiddle~40 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~40 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~30 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~30_combout ),
	.cout());
defparam \reg_no_twiddle~30 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~30 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~20 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~20_combout ),
	.cout());
defparam \reg_no_twiddle~20 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~20 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~10 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~10_combout ),
	.cout());
defparam \reg_no_twiddle~10 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~10 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~0 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~0_combout ),
	.cout());
defparam \reg_no_twiddle~0 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][0][6]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][5]~2 ),
	.combout(\reg_no_twiddle[0][0][6]~1_combout ),
	.cout(\reg_no_twiddle[0][0][6]~2 ));
defparam \reg_no_twiddle[0][0][6]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][7]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][6]~2 ),
	.combout(\reg_no_twiddle[0][0][7]~1_combout ),
	.cout(\reg_no_twiddle[0][0][7]~2 ));
defparam \reg_no_twiddle[0][0][7]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][8]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][0][7]~2 ),
	.combout(\reg_no_twiddle[0][0][8]~1_combout ),
	.cout(\reg_no_twiddle[0][0][8]~2 ));
defparam \reg_no_twiddle[0][0][8]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][0][9]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\reg_no_twiddle[0][0][8]~2 ),
	.combout(\reg_no_twiddle[0][0][9]~1_combout ),
	.cout());
defparam \reg_no_twiddle[0][0][9]~1 .lut_mask = 16'h5A5A;
defparam \reg_no_twiddle[0][0][9]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~61 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~61_combout ),
	.cout());
defparam \reg_no_twiddle~61 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~61 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~41 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~41_combout ),
	.cout());
defparam \reg_no_twiddle~41 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~41 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~31 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~31_combout ),
	.cout());
defparam \reg_no_twiddle~31 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~31 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~21 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~21_combout ),
	.cout());
defparam \reg_no_twiddle~21 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~21 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~11 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~11_combout ),
	.cout());
defparam \reg_no_twiddle~11 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~11 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][9] (
	.clk(clk),
	.d(\reg_no_twiddle~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~1 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~1_combout ),
	.cout());
defparam \reg_no_twiddle~1 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle~81 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.cin(gnd),
	.combout(\reg_no_twiddle~81_combout ),
	.cout());
defparam \reg_no_twiddle~81 .lut_mask = 16'hAAFF;
defparam \reg_no_twiddle~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][1][0]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\reg_no_twiddle~81_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\reg_no_twiddle[0][1][0]~1_combout ),
	.cout(\reg_no_twiddle[0][1][0]~2 ));
defparam \reg_no_twiddle[0][1][0]~1 .lut_mask = 16'h66EE;
defparam \reg_no_twiddle[0][1][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][1][1]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][0]~2 ),
	.combout(\reg_no_twiddle[0][1][1]~1_combout ),
	.cout(\reg_no_twiddle[0][1][1]~2 ));
defparam \reg_no_twiddle[0][1][1]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][1]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][2]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][1]~2 ),
	.combout(\reg_no_twiddle[0][1][2]~1_combout ),
	.cout(\reg_no_twiddle[0][1][2]~2 ));
defparam \reg_no_twiddle[0][1][2]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][2]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][3]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][2]~2 ),
	.combout(\reg_no_twiddle[0][1][3]~1_combout ),
	.cout(\reg_no_twiddle[0][1][3]~2 ));
defparam \reg_no_twiddle[0][1][3]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][3]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][4]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][3]~2 ),
	.combout(\reg_no_twiddle[0][1][4]~1_combout ),
	.cout(\reg_no_twiddle[0][1][4]~2 ));
defparam \reg_no_twiddle[0][1][4]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][4]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][5]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][4]~2 ),
	.combout(\reg_no_twiddle[0][1][5]~1_combout ),
	.cout(\reg_no_twiddle[0][1][5]~2 ));
defparam \reg_no_twiddle[0][1][5]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][5]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~62 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~62_combout ),
	.cout());
defparam \reg_no_twiddle~62 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~62 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~42 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~42_combout ),
	.cout());
defparam \reg_no_twiddle~42 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~42 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~32 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~32_combout ),
	.cout());
defparam \reg_no_twiddle~32 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~32 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~22 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~22_combout ),
	.cout());
defparam \reg_no_twiddle~22 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~22 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~12 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~12_combout ),
	.cout());
defparam \reg_no_twiddle~12 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~12 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][5] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~2 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~2_combout ),
	.cout());
defparam \reg_no_twiddle~2 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \reg_no_twiddle[0][1][6]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][5]~2 ),
	.combout(\reg_no_twiddle[0][1][6]~1_combout ),
	.cout(\reg_no_twiddle[0][1][6]~2 ));
defparam \reg_no_twiddle[0][1][6]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][7]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][6]~2 ),
	.combout(\reg_no_twiddle[0][1][7]~1_combout ),
	.cout(\reg_no_twiddle[0][1][7]~2 ));
defparam \reg_no_twiddle[0][1][7]~1 .lut_mask = 16'h5A5F;
defparam \reg_no_twiddle[0][1][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][8]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\reg_no_twiddle[0][1][7]~2 ),
	.combout(\reg_no_twiddle[0][1][8]~1_combout ),
	.cout(\reg_no_twiddle[0][1][8]~2 ));
defparam \reg_no_twiddle[0][1][8]~1 .lut_mask = 16'h5AAF;
defparam \reg_no_twiddle[0][1][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \reg_no_twiddle[0][1][9]~1 (
	.dataa(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\reg_no_twiddle[0][1][8]~2 ),
	.combout(\reg_no_twiddle[0][1][9]~1_combout ),
	.cout());
defparam \reg_no_twiddle[0][1][9]~1 .lut_mask = 16'h5A5A;
defparam \reg_no_twiddle[0][1][9]~1 .sum_lutc_input = "cin";

dffeas \reg_no_twiddle[0][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~63 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~63_combout ),
	.cout());
defparam \reg_no_twiddle~63 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~63 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~43 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~43_combout ),
	.cout());
defparam \reg_no_twiddle~43 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~43 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~33 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~33_combout ),
	.cout());
defparam \reg_no_twiddle~33 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~33 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~23 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~23_combout ),
	.cout());
defparam \reg_no_twiddle~23 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~23 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~13 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~13_combout ),
	.cout());
defparam \reg_no_twiddle~13 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~13 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][9] (
	.clk(clk),
	.d(\reg_no_twiddle~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][9]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][9] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][9] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~3 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~3_combout ),
	.cout());
defparam \reg_no_twiddle~3 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~3 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~64 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~64_combout ),
	.cout());
defparam \reg_no_twiddle~64 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~64 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~44 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~44_combout ),
	.cout());
defparam \reg_no_twiddle~44 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~44 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~34 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~34_combout ),
	.cout());
defparam \reg_no_twiddle~34 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~34 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~24 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~24_combout ),
	.cout());
defparam \reg_no_twiddle~24 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~24 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~14 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~14_combout ),
	.cout());
defparam \reg_no_twiddle~14 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~14 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~4 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~4_combout ),
	.cout());
defparam \reg_no_twiddle~4 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~4 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~65 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~65_combout ),
	.cout());
defparam \reg_no_twiddle~65 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~65 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~45 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~45_combout ),
	.cout());
defparam \reg_no_twiddle~45 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~45 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~35 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~35_combout ),
	.cout());
defparam \reg_no_twiddle~35 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~35 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~25 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~25_combout ),
	.cout());
defparam \reg_no_twiddle~25 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~25 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~15 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~15_combout ),
	.cout());
defparam \reg_no_twiddle~15 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~15 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][6] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~5 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~5_combout ),
	.cout());
defparam \reg_no_twiddle~5 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~5 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~66 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~66_combout ),
	.cout());
defparam \reg_no_twiddle~66 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~66 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~46 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~46_combout ),
	.cout());
defparam \reg_no_twiddle~46 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~46 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~36 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~36_combout ),
	.cout());
defparam \reg_no_twiddle~36 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~36 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~26 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~26_combout ),
	.cout());
defparam \reg_no_twiddle~26 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~26 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~16 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~16_combout ),
	.cout());
defparam \reg_no_twiddle~16 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~16 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~6 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~6_combout ),
	.cout());
defparam \reg_no_twiddle~6 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~6 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~67 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~67_combout ),
	.cout());
defparam \reg_no_twiddle~67 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~67 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~47 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~47_combout ),
	.cout());
defparam \reg_no_twiddle~47 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~47 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~37 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~37_combout ),
	.cout());
defparam \reg_no_twiddle~37 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~37 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~27 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~27_combout ),
	.cout());
defparam \reg_no_twiddle~27 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~27 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~17 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~17_combout ),
	.cout());
defparam \reg_no_twiddle~17 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~17 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][7] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~7 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~7_combout ),
	.cout());
defparam \reg_no_twiddle~7 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~7 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~68 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~68_combout ),
	.cout());
defparam \reg_no_twiddle~68 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~68 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~48 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~48_combout ),
	.cout());
defparam \reg_no_twiddle~48 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~48 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~38 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~38_combout ),
	.cout());
defparam \reg_no_twiddle~38 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~38 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~28 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~28_combout ),
	.cout());
defparam \reg_no_twiddle~28 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~28 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~18 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~18_combout ),
	.cout());
defparam \reg_no_twiddle~18 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~18 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][8] (
	.clk(clk),
	.d(\reg_no_twiddle~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~8 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~8_combout ),
	.cout());
defparam \reg_no_twiddle~8 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~8 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~69 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~69_combout ),
	.cout());
defparam \reg_no_twiddle~69 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~69 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~49 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~49_combout ),
	.cout());
defparam \reg_no_twiddle~49 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~49 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~39 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~39_combout ),
	.cout());
defparam \reg_no_twiddle~39 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~39 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~29 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~29_combout ),
	.cout());
defparam \reg_no_twiddle~29 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~29 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~19 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~19_combout ),
	.cout());
defparam \reg_no_twiddle~19 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~19 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][8] (
	.clk(clk),
	.d(\reg_no_twiddle~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][8]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][8] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][8] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~9 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~9_combout ),
	.cout());
defparam \reg_no_twiddle~9 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~9 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~112 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~112_combout ),
	.cout());
defparam \reg_no_twiddle~112 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~112 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~112_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~102 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~102_combout ),
	.cout());
defparam \reg_no_twiddle~102 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~102 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~102_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~92 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~92_combout ),
	.cout());
defparam \reg_no_twiddle~92 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~92 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~92_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~82 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~82_combout ),
	.cout());
defparam \reg_no_twiddle~82 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~82 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~70 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~70_combout ),
	.cout());
defparam \reg_no_twiddle~70 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~70 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~50 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~50_combout ),
	.cout());
defparam \reg_no_twiddle~50 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~50 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~113 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~113_combout ),
	.cout());
defparam \reg_no_twiddle~113 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~113 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~113_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~103 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~103_combout ),
	.cout());
defparam \reg_no_twiddle~103 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~103 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~103_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~93 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~93_combout ),
	.cout());
defparam \reg_no_twiddle~93 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~93 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~83 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~83_combout ),
	.cout());
defparam \reg_no_twiddle~83 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~83 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~71 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~71_combout ),
	.cout());
defparam \reg_no_twiddle~71 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~71 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][2] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~51 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~51_combout ),
	.cout());
defparam \reg_no_twiddle~51 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~51 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~114 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~114_combout ),
	.cout());
defparam \reg_no_twiddle~114 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~114 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~114_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~104 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~104_combout ),
	.cout());
defparam \reg_no_twiddle~104 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~104 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~104_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~94 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~94_combout ),
	.cout());
defparam \reg_no_twiddle~94 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~94 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~94_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~84 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~84_combout ),
	.cout());
defparam \reg_no_twiddle~84 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~84 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~72 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~72_combout ),
	.cout());
defparam \reg_no_twiddle~72 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~72 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~52 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~52_combout ),
	.cout());
defparam \reg_no_twiddle~52 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~52 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~115 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~115_combout ),
	.cout());
defparam \reg_no_twiddle~115 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~115 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~115_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~105 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~105_combout ),
	.cout());
defparam \reg_no_twiddle~105 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~105 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~105_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~95 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~95_combout ),
	.cout());
defparam \reg_no_twiddle~95 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~95 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~95_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~85 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~85_combout ),
	.cout());
defparam \reg_no_twiddle~85 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~85 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~73 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~73_combout ),
	.cout());
defparam \reg_no_twiddle~73 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~73 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][1] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~53 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~53_combout ),
	.cout());
defparam \reg_no_twiddle~53 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~53 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~116 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~116_combout ),
	.cout());
defparam \reg_no_twiddle~116 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~116 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~116_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~106 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~106_combout ),
	.cout());
defparam \reg_no_twiddle~106 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~106 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~106_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~96 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~96_combout ),
	.cout());
defparam \reg_no_twiddle~96 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~96 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~86 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~86_combout ),
	.cout());
defparam \reg_no_twiddle~86 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~86 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~74 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~74_combout ),
	.cout());
defparam \reg_no_twiddle~74 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~74 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~54 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~54_combout ),
	.cout());
defparam \reg_no_twiddle~54 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~54 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~117 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~117_combout ),
	.cout());
defparam \reg_no_twiddle~117 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~117 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~117_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~107 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~107_combout ),
	.cout());
defparam \reg_no_twiddle~107 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~107 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~107_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~97 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~97_combout ),
	.cout());
defparam \reg_no_twiddle~97 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~97 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~97_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~87 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~87_combout ),
	.cout());
defparam \reg_no_twiddle~87 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~87 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~75 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~75_combout ),
	.cout());
defparam \reg_no_twiddle~75 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~75 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][0] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~55 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~55_combout ),
	.cout());
defparam \reg_no_twiddle~55 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~55 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~118 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~118_combout ),
	.cout());
defparam \reg_no_twiddle~118 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~118 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~118_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~108 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~108_combout ),
	.cout());
defparam \reg_no_twiddle~108 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~108 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~108_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~98 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~98_combout ),
	.cout());
defparam \reg_no_twiddle~98 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~98 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~98_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~88 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~88_combout ),
	.cout());
defparam \reg_no_twiddle~88 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~88 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~76 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~76_combout ),
	.cout());
defparam \reg_no_twiddle~76 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~76 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~56 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~56_combout ),
	.cout());
defparam \reg_no_twiddle~56 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~56 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~119 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~119_combout ),
	.cout());
defparam \reg_no_twiddle~119 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~119 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~119_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~109 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~109_combout ),
	.cout());
defparam \reg_no_twiddle~109 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~109 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~109_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~99 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~99_combout ),
	.cout());
defparam \reg_no_twiddle~99 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~99 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~99_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~89 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~89_combout ),
	.cout());
defparam \reg_no_twiddle~89 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~89 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~89_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~77 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~77_combout ),
	.cout());
defparam \reg_no_twiddle~77 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~77 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][4] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~57 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~57_combout ),
	.cout());
defparam \reg_no_twiddle~57 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~57 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~120 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~120_combout ),
	.cout());
defparam \reg_no_twiddle~120 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~120 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~120_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~110 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~110_combout ),
	.cout());
defparam \reg_no_twiddle~110 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~110 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~110_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~100 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~100_combout ),
	.cout());
defparam \reg_no_twiddle~100 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~100 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~100_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~90 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~90_combout ),
	.cout());
defparam \reg_no_twiddle~90 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~90 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~78 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~78_combout ),
	.cout());
defparam \reg_no_twiddle~78 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~78 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~58 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~58_combout ),
	.cout());
defparam \reg_no_twiddle~58 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~58 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[0][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[0][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~121 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[0][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~121_combout ),
	.cout());
defparam \reg_no_twiddle~121 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~121 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[1][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~121_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[1][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~111 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[1][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~111_combout ),
	.cout());
defparam \reg_no_twiddle~111 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~111 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[2][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~111_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[2][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~101 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[2][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~101_combout ),
	.cout());
defparam \reg_no_twiddle~101 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~101 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[3][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[3][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~91 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[3][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~91_combout ),
	.cout());
defparam \reg_no_twiddle~91 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~91 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[4][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~91_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[4][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~79 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[4][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~79_combout ),
	.cout());
defparam \reg_no_twiddle~79 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~79 .sum_lutc_input = "datac";

dffeas \reg_no_twiddle[5][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\reg_no_twiddle[5][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][3] .power_up = "low";

cycloneive_lcell_comb \reg_no_twiddle~59 (
	.dataa(reset_n),
	.datab(\reg_no_twiddle[5][1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_no_twiddle~59_combout ),
	.cout());
defparam \reg_no_twiddle~59 .lut_mask = 16'hEEEE;
defparam \reg_no_twiddle~59 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_bfp_i (
	r_array_out_7_2,
	r_array_out_7_0,
	r_array_out_6_2,
	r_array_out_6_0,
	r_array_out_5_2,
	r_array_out_5_0,
	r_array_out_4_2,
	r_array_out_4_0,
	r_array_out_3_2,
	r_array_out_3_0,
	r_array_out_2_2,
	r_array_out_2_0,
	r_array_out_7_3,
	r_array_out_7_1,
	r_array_out_6_3,
	r_array_out_6_1,
	r_array_out_5_3,
	r_array_out_5_1,
	r_array_out_4_3,
	r_array_out_4_1,
	r_array_out_3_3,
	r_array_out_3_1,
	r_array_out_2_3,
	r_array_out_2_1,
	i_array_out_7_2,
	i_array_out_7_0,
	i_array_out_6_2,
	i_array_out_6_0,
	i_array_out_5_2,
	i_array_out_5_0,
	i_array_out_4_2,
	i_array_out_4_0,
	i_array_out_3_2,
	i_array_out_3_0,
	i_array_out_2_2,
	i_array_out_2_0,
	i_array_out_7_3,
	i_array_out_7_1,
	i_array_out_6_3,
	i_array_out_6_1,
	i_array_out_5_3,
	i_array_out_5_1,
	i_array_out_4_3,
	i_array_out_4_1,
	i_array_out_3_3,
	i_array_out_3_1,
	i_array_out_2_3,
	i_array_out_2_1,
	ram_in_reg_7_0,
	ram_in_reg_5_0,
	ram_in_reg_6_0,
	ram_in_reg_8_0,
	ram_in_reg_4_0,
	ram_in_reg_7_2,
	ram_in_reg_5_2,
	ram_in_reg_6_2,
	ram_in_reg_8_2,
	ram_in_reg_4_2,
	ram_in_reg_3_2,
	ram_in_reg_3_0,
	ram_in_reg_2_2,
	ram_in_reg_2_0,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	ram_in_reg_0_2,
	ram_in_reg_0_0,
	ram_in_reg_7_1,
	ram_in_reg_5_1,
	ram_in_reg_6_1,
	ram_in_reg_8_1,
	ram_in_reg_4_1,
	ram_in_reg_7_3,
	ram_in_reg_5_3,
	ram_in_reg_6_3,
	ram_in_reg_8_3,
	ram_in_reg_4_3,
	ram_in_reg_3_3,
	ram_in_reg_3_1,
	ram_in_reg_2_3,
	ram_in_reg_2_1,
	ram_in_reg_1_3,
	ram_in_reg_1_1,
	ram_in_reg_0_3,
	ram_in_reg_0_1,
	ram_in_reg_9_0,
	ram_in_reg_9_2,
	ram_in_reg_9_1,
	ram_in_reg_9_3,
	ram_in_reg_5_4,
	ram_in_reg_6_4,
	ram_in_reg_7_4,
	ram_in_reg_8_4,
	ram_in_reg_4_4,
	ram_in_reg_5_6,
	ram_in_reg_6_6,
	ram_in_reg_7_6,
	ram_in_reg_8_6,
	ram_in_reg_4_6,
	ram_in_reg_3_6,
	ram_in_reg_3_4,
	ram_in_reg_2_6,
	ram_in_reg_2_4,
	ram_in_reg_1_6,
	ram_in_reg_1_4,
	ram_in_reg_0_6,
	ram_in_reg_0_4,
	ram_in_reg_5_5,
	ram_in_reg_6_5,
	ram_in_reg_7_5,
	ram_in_reg_8_5,
	ram_in_reg_4_5,
	ram_in_reg_5_7,
	ram_in_reg_6_7,
	ram_in_reg_7_7,
	ram_in_reg_8_7,
	ram_in_reg_4_7,
	ram_in_reg_3_7,
	ram_in_reg_3_5,
	ram_in_reg_2_7,
	ram_in_reg_2_5,
	ram_in_reg_1_7,
	ram_in_reg_1_5,
	ram_in_reg_0_7,
	ram_in_reg_0_5,
	ram_in_reg_9_4,
	ram_in_reg_9_6,
	ram_in_reg_9_5,
	ram_in_reg_9_7,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	r_array_out_8_0,
	r_array_out_8_2,
	r_array_out_1_0,
	r_array_out_1_2,
	r_array_out_0_0,
	r_array_out_0_2,
	r_array_out_8_1,
	r_array_out_8_3,
	r_array_out_1_1,
	r_array_out_1_3,
	r_array_out_0_1,
	r_array_out_0_3,
	r_array_out_9_0,
	r_array_out_9_2,
	r_array_out_9_1,
	r_array_out_9_3,
	i_array_out_8_0,
	i_array_out_8_2,
	i_array_out_1_0,
	i_array_out_1_2,
	i_array_out_0_0,
	i_array_out_0_2,
	i_array_out_8_1,
	i_array_out_8_3,
	i_array_out_1_1,
	i_array_out_1_3,
	i_array_out_0_1,
	i_array_out_0_3,
	i_array_out_9_0,
	i_array_out_9_2,
	i_array_out_9_1,
	i_array_out_9_3,
	clk)/* synthesis synthesis_greybox=1 */;
output 	r_array_out_7_2;
output 	r_array_out_7_0;
output 	r_array_out_6_2;
output 	r_array_out_6_0;
output 	r_array_out_5_2;
output 	r_array_out_5_0;
output 	r_array_out_4_2;
output 	r_array_out_4_0;
output 	r_array_out_3_2;
output 	r_array_out_3_0;
output 	r_array_out_2_2;
output 	r_array_out_2_0;
output 	r_array_out_7_3;
output 	r_array_out_7_1;
output 	r_array_out_6_3;
output 	r_array_out_6_1;
output 	r_array_out_5_3;
output 	r_array_out_5_1;
output 	r_array_out_4_3;
output 	r_array_out_4_1;
output 	r_array_out_3_3;
output 	r_array_out_3_1;
output 	r_array_out_2_3;
output 	r_array_out_2_1;
output 	i_array_out_7_2;
output 	i_array_out_7_0;
output 	i_array_out_6_2;
output 	i_array_out_6_0;
output 	i_array_out_5_2;
output 	i_array_out_5_0;
output 	i_array_out_4_2;
output 	i_array_out_4_0;
output 	i_array_out_3_2;
output 	i_array_out_3_0;
output 	i_array_out_2_2;
output 	i_array_out_2_0;
output 	i_array_out_7_3;
output 	i_array_out_7_1;
output 	i_array_out_6_3;
output 	i_array_out_6_1;
output 	i_array_out_5_3;
output 	i_array_out_5_1;
output 	i_array_out_4_3;
output 	i_array_out_4_1;
output 	i_array_out_3_3;
output 	i_array_out_3_1;
output 	i_array_out_2_3;
output 	i_array_out_2_1;
input 	ram_in_reg_7_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_6_0;
input 	ram_in_reg_8_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_6_2;
input 	ram_in_reg_8_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_2_0;
input 	ram_in_reg_1_2;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_6_1;
input 	ram_in_reg_8_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_6_3;
input 	ram_in_reg_8_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_1;
input 	ram_in_reg_2_3;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_9_0;
input 	ram_in_reg_9_2;
input 	ram_in_reg_9_1;
input 	ram_in_reg_9_3;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_4;
input 	ram_in_reg_8_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_6;
input 	ram_in_reg_8_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_3_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_2_4;
input 	ram_in_reg_1_6;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_5;
input 	ram_in_reg_8_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_7;
input 	ram_in_reg_8_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_5;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_9_4;
input 	ram_in_reg_9_6;
input 	ram_in_reg_9_5;
input 	ram_in_reg_9_7;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	r_array_out_8_0;
output 	r_array_out_8_2;
output 	r_array_out_1_0;
output 	r_array_out_1_2;
output 	r_array_out_0_0;
output 	r_array_out_0_2;
output 	r_array_out_8_1;
output 	r_array_out_8_3;
output 	r_array_out_1_1;
output 	r_array_out_1_3;
output 	r_array_out_0_1;
output 	r_array_out_0_3;
output 	r_array_out_9_0;
output 	r_array_out_9_2;
output 	r_array_out_9_1;
output 	r_array_out_9_3;
output 	i_array_out_8_0;
output 	i_array_out_8_2;
output 	i_array_out_1_0;
output 	i_array_out_1_2;
output 	i_array_out_0_0;
output 	i_array_out_0_2;
output 	i_array_out_8_1;
output 	i_array_out_8_3;
output 	i_array_out_1_1;
output 	i_array_out_1_3;
output 	i_array_out_0_1;
output 	i_array_out_0_3;
output 	i_array_out_9_0;
output 	i_array_out_9_2;
output 	i_array_out_9_1;
output 	i_array_out_9_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux22~0_combout ;
wire \Mux20~1_combout ;
wire \Mux22~1_combout ;
wire \Mux2~0_combout ;
wire \Mux0~1_combout ;
wire \Mux2~1_combout ;
wire \Mux23~0_combout ;
wire \Mux20~0_combout ;
wire \Mux23~1_combout ;
wire \Mux3~0_combout ;
wire \Mux0~0_combout ;
wire \Mux3~1_combout ;
wire \Mux24~0_combout ;
wire \Mux25~0_combout ;
wire \Mux24~1_combout ;
wire \Mux4~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~1_combout ;
wire \Mux26~0_combout ;
wire \Mux25~1_combout ;
wire \Mux6~0_combout ;
wire \Mux5~1_combout ;
wire \Mux26~1_combout ;
wire \Mux26~2_combout ;
wire \Mux6~1_combout ;
wire \Mux6~2_combout ;
wire \Mux27~0_combout ;
wire \Mux7~0_combout ;
wire \Mux32~0_combout ;
wire \Mux30~1_combout ;
wire \Mux32~1_combout ;
wire \Mux12~0_combout ;
wire \Mux10~1_combout ;
wire \Mux12~1_combout ;
wire \Mux33~0_combout ;
wire \Mux30~0_combout ;
wire \Mux33~1_combout ;
wire \Mux13~0_combout ;
wire \Mux10~0_combout ;
wire \Mux13~1_combout ;
wire \Mux34~0_combout ;
wire \Mux35~0_combout ;
wire \Mux34~1_combout ;
wire \Mux14~0_combout ;
wire \Mux15~0_combout ;
wire \Mux14~1_combout ;
wire \Mux36~0_combout ;
wire \Mux35~1_combout ;
wire \Mux16~0_combout ;
wire \Mux15~1_combout ;
wire \Mux36~1_combout ;
wire \Mux36~2_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \Mux37~0_combout ;
wire \Mux17~0_combout ;
wire \Mux62~0_combout ;
wire \Mux60~1_combout ;
wire \Mux62~1_combout ;
wire \Mux42~0_combout ;
wire \Mux40~1_combout ;
wire \Mux42~1_combout ;
wire \Mux63~0_combout ;
wire \Mux60~0_combout ;
wire \Mux63~1_combout ;
wire \Mux43~0_combout ;
wire \Mux40~0_combout ;
wire \Mux43~1_combout ;
wire \Mux64~0_combout ;
wire \Mux65~0_combout ;
wire \Mux64~1_combout ;
wire \Mux44~0_combout ;
wire \Mux45~0_combout ;
wire \Mux44~1_combout ;
wire \Mux66~0_combout ;
wire \Mux65~1_combout ;
wire \Mux46~0_combout ;
wire \Mux45~1_combout ;
wire \Mux66~1_combout ;
wire \Mux66~2_combout ;
wire \Mux46~1_combout ;
wire \Mux46~2_combout ;
wire \Mux67~0_combout ;
wire \Mux47~0_combout ;
wire \Mux72~0_combout ;
wire \Mux70~1_combout ;
wire \Mux72~1_combout ;
wire \Mux52~0_combout ;
wire \Mux50~1_combout ;
wire \Mux52~1_combout ;
wire \Mux73~0_combout ;
wire \Mux70~0_combout ;
wire \Mux73~1_combout ;
wire \Mux53~0_combout ;
wire \Mux50~0_combout ;
wire \Mux53~1_combout ;
wire \Mux74~0_combout ;
wire \Mux75~0_combout ;
wire \Mux74~1_combout ;
wire \Mux54~0_combout ;
wire \Mux55~0_combout ;
wire \Mux54~1_combout ;
wire \Mux76~0_combout ;
wire \Mux75~1_combout ;
wire \Mux56~0_combout ;
wire \Mux55~1_combout ;
wire \Mux76~1_combout ;
wire \Mux76~2_combout ;
wire \Mux56~1_combout ;
wire \Mux56~2_combout ;
wire \Mux77~0_combout ;
wire \Mux57~0_combout ;
wire \i_array_out[2][9]~0_combout ;
wire \i_array_out[2][9]~1_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux8~0_combout ;
wire \Mux28~0_combout ;
wire \Mux9~0_combout ;
wire \Mux29~0_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux18~0_combout ;
wire \Mux38~0_combout ;
wire \Mux19~0_combout ;
wire \Mux39~0_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux48~0_combout ;
wire \Mux68~0_combout ;
wire \Mux49~0_combout ;
wire \Mux69~0_combout ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \Mux71~0_combout ;
wire \Mux71~1_combout ;
wire \Mux58~0_combout ;
wire \Mux78~0_combout ;
wire \Mux59~0_combout ;
wire \Mux79~0_combout ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \Mux70~2_combout ;
wire \Mux70~3_combout ;


dffeas \r_array_out[2][7] (
	.clk(clk),
	.d(\Mux22~1_combout ),
	.asdata(ram_in_reg_3_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_7_2),
	.prn(vcc));
defparam \r_array_out[2][7] .is_wysiwyg = "true";
defparam \r_array_out[2][7] .power_up = "low";

dffeas \r_array_out[0][7] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(ram_in_reg_3_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_7_0),
	.prn(vcc));
defparam \r_array_out[0][7] .is_wysiwyg = "true";
defparam \r_array_out[0][7] .power_up = "low";

dffeas \r_array_out[2][6] (
	.clk(clk),
	.d(\Mux23~1_combout ),
	.asdata(ram_in_reg_2_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_6_2),
	.prn(vcc));
defparam \r_array_out[2][6] .is_wysiwyg = "true";
defparam \r_array_out[2][6] .power_up = "low";

dffeas \r_array_out[0][6] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(ram_in_reg_2_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_6_0),
	.prn(vcc));
defparam \r_array_out[0][6] .is_wysiwyg = "true";
defparam \r_array_out[0][6] .power_up = "low";

dffeas \r_array_out[2][5] (
	.clk(clk),
	.d(\Mux24~1_combout ),
	.asdata(ram_in_reg_1_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_2),
	.prn(vcc));
defparam \r_array_out[2][5] .is_wysiwyg = "true";
defparam \r_array_out[2][5] .power_up = "low";

dffeas \r_array_out[0][5] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(ram_in_reg_1_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_0),
	.prn(vcc));
defparam \r_array_out[0][5] .is_wysiwyg = "true";
defparam \r_array_out[0][5] .power_up = "low";

dffeas \r_array_out[2][4] (
	.clk(clk),
	.d(\Mux25~1_combout ),
	.asdata(ram_in_reg_0_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_2),
	.prn(vcc));
defparam \r_array_out[2][4] .is_wysiwyg = "true";
defparam \r_array_out[2][4] .power_up = "low";

dffeas \r_array_out[0][4] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(ram_in_reg_0_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_0),
	.prn(vcc));
defparam \r_array_out[0][4] .is_wysiwyg = "true";
defparam \r_array_out[0][4] .power_up = "low";

dffeas \r_array_out[2][3] (
	.clk(clk),
	.d(\Mux26~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_3_2),
	.prn(vcc));
defparam \r_array_out[2][3] .is_wysiwyg = "true";
defparam \r_array_out[2][3] .power_up = "low";

dffeas \r_array_out[0][3] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_3_0),
	.prn(vcc));
defparam \r_array_out[0][3] .is_wysiwyg = "true";
defparam \r_array_out[0][3] .power_up = "low";

dffeas \r_array_out[2][2] (
	.clk(clk),
	.d(\Mux27~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_2_2),
	.prn(vcc));
defparam \r_array_out[2][2] .is_wysiwyg = "true";
defparam \r_array_out[2][2] .power_up = "low";

dffeas \r_array_out[0][2] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_2_0),
	.prn(vcc));
defparam \r_array_out[0][2] .is_wysiwyg = "true";
defparam \r_array_out[0][2] .power_up = "low";

dffeas \r_array_out[3][7] (
	.clk(clk),
	.d(\Mux32~1_combout ),
	.asdata(ram_in_reg_3_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_7_3),
	.prn(vcc));
defparam \r_array_out[3][7] .is_wysiwyg = "true";
defparam \r_array_out[3][7] .power_up = "low";

dffeas \r_array_out[1][7] (
	.clk(clk),
	.d(\Mux12~1_combout ),
	.asdata(ram_in_reg_3_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_7_1),
	.prn(vcc));
defparam \r_array_out[1][7] .is_wysiwyg = "true";
defparam \r_array_out[1][7] .power_up = "low";

dffeas \r_array_out[3][6] (
	.clk(clk),
	.d(\Mux33~1_combout ),
	.asdata(ram_in_reg_2_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_6_3),
	.prn(vcc));
defparam \r_array_out[3][6] .is_wysiwyg = "true";
defparam \r_array_out[3][6] .power_up = "low";

dffeas \r_array_out[1][6] (
	.clk(clk),
	.d(\Mux13~1_combout ),
	.asdata(ram_in_reg_2_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_6_1),
	.prn(vcc));
defparam \r_array_out[1][6] .is_wysiwyg = "true";
defparam \r_array_out[1][6] .power_up = "low";

dffeas \r_array_out[3][5] (
	.clk(clk),
	.d(\Mux34~1_combout ),
	.asdata(ram_in_reg_1_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_3),
	.prn(vcc));
defparam \r_array_out[3][5] .is_wysiwyg = "true";
defparam \r_array_out[3][5] .power_up = "low";

dffeas \r_array_out[1][5] (
	.clk(clk),
	.d(\Mux14~1_combout ),
	.asdata(ram_in_reg_1_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_5_1),
	.prn(vcc));
defparam \r_array_out[1][5] .is_wysiwyg = "true";
defparam \r_array_out[1][5] .power_up = "low";

dffeas \r_array_out[3][4] (
	.clk(clk),
	.d(\Mux35~1_combout ),
	.asdata(ram_in_reg_0_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_3),
	.prn(vcc));
defparam \r_array_out[3][4] .is_wysiwyg = "true";
defparam \r_array_out[3][4] .power_up = "low";

dffeas \r_array_out[1][4] (
	.clk(clk),
	.d(\Mux15~1_combout ),
	.asdata(ram_in_reg_0_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(r_array_out_4_1),
	.prn(vcc));
defparam \r_array_out[1][4] .is_wysiwyg = "true";
defparam \r_array_out[1][4] .power_up = "low";

dffeas \r_array_out[3][3] (
	.clk(clk),
	.d(\Mux36~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_3_3),
	.prn(vcc));
defparam \r_array_out[3][3] .is_wysiwyg = "true";
defparam \r_array_out[3][3] .power_up = "low";

dffeas \r_array_out[1][3] (
	.clk(clk),
	.d(\Mux16~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_3_1),
	.prn(vcc));
defparam \r_array_out[1][3] .is_wysiwyg = "true";
defparam \r_array_out[1][3] .power_up = "low";

dffeas \r_array_out[3][2] (
	.clk(clk),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_2_3),
	.prn(vcc));
defparam \r_array_out[3][2] .is_wysiwyg = "true";
defparam \r_array_out[3][2] .power_up = "low";

dffeas \r_array_out[1][2] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_2_1),
	.prn(vcc));
defparam \r_array_out[1][2] .is_wysiwyg = "true";
defparam \r_array_out[1][2] .power_up = "low";

dffeas \i_array_out[2][7] (
	.clk(clk),
	.d(\Mux62~1_combout ),
	.asdata(ram_in_reg_3_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_7_2),
	.prn(vcc));
defparam \i_array_out[2][7] .is_wysiwyg = "true";
defparam \i_array_out[2][7] .power_up = "low";

dffeas \i_array_out[0][7] (
	.clk(clk),
	.d(\Mux42~1_combout ),
	.asdata(ram_in_reg_3_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_7_0),
	.prn(vcc));
defparam \i_array_out[0][7] .is_wysiwyg = "true";
defparam \i_array_out[0][7] .power_up = "low";

dffeas \i_array_out[2][6] (
	.clk(clk),
	.d(\Mux63~1_combout ),
	.asdata(ram_in_reg_2_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_6_2),
	.prn(vcc));
defparam \i_array_out[2][6] .is_wysiwyg = "true";
defparam \i_array_out[2][6] .power_up = "low";

dffeas \i_array_out[0][6] (
	.clk(clk),
	.d(\Mux43~1_combout ),
	.asdata(ram_in_reg_2_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_6_0),
	.prn(vcc));
defparam \i_array_out[0][6] .is_wysiwyg = "true";
defparam \i_array_out[0][6] .power_up = "low";

dffeas \i_array_out[2][5] (
	.clk(clk),
	.d(\Mux64~1_combout ),
	.asdata(ram_in_reg_1_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_2),
	.prn(vcc));
defparam \i_array_out[2][5] .is_wysiwyg = "true";
defparam \i_array_out[2][5] .power_up = "low";

dffeas \i_array_out[0][5] (
	.clk(clk),
	.d(\Mux44~1_combout ),
	.asdata(ram_in_reg_1_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_0),
	.prn(vcc));
defparam \i_array_out[0][5] .is_wysiwyg = "true";
defparam \i_array_out[0][5] .power_up = "low";

dffeas \i_array_out[2][4] (
	.clk(clk),
	.d(\Mux65~1_combout ),
	.asdata(ram_in_reg_0_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_2),
	.prn(vcc));
defparam \i_array_out[2][4] .is_wysiwyg = "true";
defparam \i_array_out[2][4] .power_up = "low";

dffeas \i_array_out[0][4] (
	.clk(clk),
	.d(\Mux45~1_combout ),
	.asdata(ram_in_reg_0_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_0),
	.prn(vcc));
defparam \i_array_out[0][4] .is_wysiwyg = "true";
defparam \i_array_out[0][4] .power_up = "low";

dffeas \i_array_out[2][3] (
	.clk(clk),
	.d(\Mux66~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_3_2),
	.prn(vcc));
defparam \i_array_out[2][3] .is_wysiwyg = "true";
defparam \i_array_out[2][3] .power_up = "low";

dffeas \i_array_out[0][3] (
	.clk(clk),
	.d(\Mux46~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_3_0),
	.prn(vcc));
defparam \i_array_out[0][3] .is_wysiwyg = "true";
defparam \i_array_out[0][3] .power_up = "low";

dffeas \i_array_out[2][2] (
	.clk(clk),
	.d(\Mux67~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_2_2),
	.prn(vcc));
defparam \i_array_out[2][2] .is_wysiwyg = "true";
defparam \i_array_out[2][2] .power_up = "low";

dffeas \i_array_out[0][2] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_2_0),
	.prn(vcc));
defparam \i_array_out[0][2] .is_wysiwyg = "true";
defparam \i_array_out[0][2] .power_up = "low";

dffeas \i_array_out[3][7] (
	.clk(clk),
	.d(\Mux72~1_combout ),
	.asdata(ram_in_reg_3_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_7_3),
	.prn(vcc));
defparam \i_array_out[3][7] .is_wysiwyg = "true";
defparam \i_array_out[3][7] .power_up = "low";

dffeas \i_array_out[1][7] (
	.clk(clk),
	.d(\Mux52~1_combout ),
	.asdata(ram_in_reg_3_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_7_1),
	.prn(vcc));
defparam \i_array_out[1][7] .is_wysiwyg = "true";
defparam \i_array_out[1][7] .power_up = "low";

dffeas \i_array_out[3][6] (
	.clk(clk),
	.d(\Mux73~1_combout ),
	.asdata(ram_in_reg_2_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_6_3),
	.prn(vcc));
defparam \i_array_out[3][6] .is_wysiwyg = "true";
defparam \i_array_out[3][6] .power_up = "low";

dffeas \i_array_out[1][6] (
	.clk(clk),
	.d(\Mux53~1_combout ),
	.asdata(ram_in_reg_2_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_6_1),
	.prn(vcc));
defparam \i_array_out[1][6] .is_wysiwyg = "true";
defparam \i_array_out[1][6] .power_up = "low";

dffeas \i_array_out[3][5] (
	.clk(clk),
	.d(\Mux74~1_combout ),
	.asdata(ram_in_reg_1_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_3),
	.prn(vcc));
defparam \i_array_out[3][5] .is_wysiwyg = "true";
defparam \i_array_out[3][5] .power_up = "low";

dffeas \i_array_out[1][5] (
	.clk(clk),
	.d(\Mux54~1_combout ),
	.asdata(ram_in_reg_1_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_5_1),
	.prn(vcc));
defparam \i_array_out[1][5] .is_wysiwyg = "true";
defparam \i_array_out[1][5] .power_up = "low";

dffeas \i_array_out[3][4] (
	.clk(clk),
	.d(\Mux75~1_combout ),
	.asdata(ram_in_reg_0_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_3),
	.prn(vcc));
defparam \i_array_out[3][4] .is_wysiwyg = "true";
defparam \i_array_out[3][4] .power_up = "low";

dffeas \i_array_out[1][4] (
	.clk(clk),
	.d(\Mux55~1_combout ),
	.asdata(ram_in_reg_0_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(global_clock_enable),
	.q(i_array_out_4_1),
	.prn(vcc));
defparam \i_array_out[1][4] .is_wysiwyg = "true";
defparam \i_array_out[1][4] .power_up = "low";

dffeas \i_array_out[3][3] (
	.clk(clk),
	.d(\Mux76~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_3_3),
	.prn(vcc));
defparam \i_array_out[3][3] .is_wysiwyg = "true";
defparam \i_array_out[3][3] .power_up = "low";

dffeas \i_array_out[1][3] (
	.clk(clk),
	.d(\Mux56~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_3_1),
	.prn(vcc));
defparam \i_array_out[1][3] .is_wysiwyg = "true";
defparam \i_array_out[1][3] .power_up = "low";

dffeas \i_array_out[3][2] (
	.clk(clk),
	.d(\Mux77~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_2_3),
	.prn(vcc));
defparam \i_array_out[3][2] .is_wysiwyg = "true";
defparam \i_array_out[3][2] .power_up = "low";

dffeas \i_array_out[1][2] (
	.clk(clk),
	.d(\Mux57~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_2_1),
	.prn(vcc));
defparam \i_array_out[1][2] .is_wysiwyg = "true";
defparam \i_array_out[1][2] .power_up = "low";

dffeas \r_array_out[0][8] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_8_0),
	.prn(vcc));
defparam \r_array_out[0][8] .is_wysiwyg = "true";
defparam \r_array_out[0][8] .power_up = "low";

dffeas \r_array_out[2][8] (
	.clk(clk),
	.d(\Mux21~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_8_2),
	.prn(vcc));
defparam \r_array_out[2][8] .is_wysiwyg = "true";
defparam \r_array_out[2][8] .power_up = "low";

dffeas \r_array_out[0][1] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_0),
	.prn(vcc));
defparam \r_array_out[0][1] .is_wysiwyg = "true";
defparam \r_array_out[0][1] .power_up = "low";

dffeas \r_array_out[2][1] (
	.clk(clk),
	.d(\Mux28~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_2),
	.prn(vcc));
defparam \r_array_out[2][1] .is_wysiwyg = "true";
defparam \r_array_out[2][1] .power_up = "low";

dffeas \r_array_out[0][0] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_0),
	.prn(vcc));
defparam \r_array_out[0][0] .is_wysiwyg = "true";
defparam \r_array_out[0][0] .power_up = "low";

dffeas \r_array_out[2][0] (
	.clk(clk),
	.d(\Mux29~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_2),
	.prn(vcc));
defparam \r_array_out[2][0] .is_wysiwyg = "true";
defparam \r_array_out[2][0] .power_up = "low";

dffeas \r_array_out[1][8] (
	.clk(clk),
	.d(\Mux11~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_8_1),
	.prn(vcc));
defparam \r_array_out[1][8] .is_wysiwyg = "true";
defparam \r_array_out[1][8] .power_up = "low";

dffeas \r_array_out[3][8] (
	.clk(clk),
	.d(\Mux31~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_8_3),
	.prn(vcc));
defparam \r_array_out[3][8] .is_wysiwyg = "true";
defparam \r_array_out[3][8] .power_up = "low";

dffeas \r_array_out[1][1] (
	.clk(clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_1),
	.prn(vcc));
defparam \r_array_out[1][1] .is_wysiwyg = "true";
defparam \r_array_out[1][1] .power_up = "low";

dffeas \r_array_out[3][1] (
	.clk(clk),
	.d(\Mux38~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_1_3),
	.prn(vcc));
defparam \r_array_out[3][1] .is_wysiwyg = "true";
defparam \r_array_out[3][1] .power_up = "low";

dffeas \r_array_out[1][0] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_1),
	.prn(vcc));
defparam \r_array_out[1][0] .is_wysiwyg = "true";
defparam \r_array_out[1][0] .power_up = "low";

dffeas \r_array_out[3][0] (
	.clk(clk),
	.d(\Mux39~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_0_3),
	.prn(vcc));
defparam \r_array_out[3][0] .is_wysiwyg = "true";
defparam \r_array_out[3][0] .power_up = "low";

dffeas \r_array_out[0][9] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_9_0),
	.prn(vcc));
defparam \r_array_out[0][9] .is_wysiwyg = "true";
defparam \r_array_out[0][9] .power_up = "low";

dffeas \r_array_out[2][9] (
	.clk(clk),
	.d(\Mux20~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_9_2),
	.prn(vcc));
defparam \r_array_out[2][9] .is_wysiwyg = "true";
defparam \r_array_out[2][9] .power_up = "low";

dffeas \r_array_out[1][9] (
	.clk(clk),
	.d(\Mux10~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_9_1),
	.prn(vcc));
defparam \r_array_out[1][9] .is_wysiwyg = "true";
defparam \r_array_out[1][9] .power_up = "low";

dffeas \r_array_out[3][9] (
	.clk(clk),
	.d(\Mux30~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(r_array_out_9_3),
	.prn(vcc));
defparam \r_array_out[3][9] .is_wysiwyg = "true";
defparam \r_array_out[3][9] .power_up = "low";

dffeas \i_array_out[0][8] (
	.clk(clk),
	.d(\Mux41~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_8_0),
	.prn(vcc));
defparam \i_array_out[0][8] .is_wysiwyg = "true";
defparam \i_array_out[0][8] .power_up = "low";

dffeas \i_array_out[2][8] (
	.clk(clk),
	.d(\Mux61~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_8_2),
	.prn(vcc));
defparam \i_array_out[2][8] .is_wysiwyg = "true";
defparam \i_array_out[2][8] .power_up = "low";

dffeas \i_array_out[0][1] (
	.clk(clk),
	.d(\Mux48~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_0),
	.prn(vcc));
defparam \i_array_out[0][1] .is_wysiwyg = "true";
defparam \i_array_out[0][1] .power_up = "low";

dffeas \i_array_out[2][1] (
	.clk(clk),
	.d(\Mux68~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_2),
	.prn(vcc));
defparam \i_array_out[2][1] .is_wysiwyg = "true";
defparam \i_array_out[2][1] .power_up = "low";

dffeas \i_array_out[0][0] (
	.clk(clk),
	.d(\Mux49~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_0),
	.prn(vcc));
defparam \i_array_out[0][0] .is_wysiwyg = "true";
defparam \i_array_out[0][0] .power_up = "low";

dffeas \i_array_out[2][0] (
	.clk(clk),
	.d(\Mux69~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_2),
	.prn(vcc));
defparam \i_array_out[2][0] .is_wysiwyg = "true";
defparam \i_array_out[2][0] .power_up = "low";

dffeas \i_array_out[1][8] (
	.clk(clk),
	.d(\Mux51~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_8_1),
	.prn(vcc));
defparam \i_array_out[1][8] .is_wysiwyg = "true";
defparam \i_array_out[1][8] .power_up = "low";

dffeas \i_array_out[3][8] (
	.clk(clk),
	.d(\Mux71~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_8_3),
	.prn(vcc));
defparam \i_array_out[3][8] .is_wysiwyg = "true";
defparam \i_array_out[3][8] .power_up = "low";

dffeas \i_array_out[1][1] (
	.clk(clk),
	.d(\Mux58~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_1),
	.prn(vcc));
defparam \i_array_out[1][1] .is_wysiwyg = "true";
defparam \i_array_out[1][1] .power_up = "low";

dffeas \i_array_out[3][1] (
	.clk(clk),
	.d(\Mux78~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_1_3),
	.prn(vcc));
defparam \i_array_out[3][1] .is_wysiwyg = "true";
defparam \i_array_out[3][1] .power_up = "low";

dffeas \i_array_out[1][0] (
	.clk(clk),
	.d(\Mux59~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_1),
	.prn(vcc));
defparam \i_array_out[1][0] .is_wysiwyg = "true";
defparam \i_array_out[1][0] .power_up = "low";

dffeas \i_array_out[3][0] (
	.clk(clk),
	.d(\Mux79~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_0_3),
	.prn(vcc));
defparam \i_array_out[3][0] .is_wysiwyg = "true";
defparam \i_array_out[3][0] .power_up = "low";

dffeas \i_array_out[0][9] (
	.clk(clk),
	.d(\Mux40~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_9_0),
	.prn(vcc));
defparam \i_array_out[0][9] .is_wysiwyg = "true";
defparam \i_array_out[0][9] .power_up = "low";

dffeas \i_array_out[2][9] (
	.clk(clk),
	.d(\Mux60~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_9_2),
	.prn(vcc));
defparam \i_array_out[2][9] .is_wysiwyg = "true";
defparam \i_array_out[2][9] .power_up = "low";

dffeas \i_array_out[1][9] (
	.clk(clk),
	.d(\Mux50~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_9_1),
	.prn(vcc));
defparam \i_array_out[1][9] .is_wysiwyg = "true";
defparam \i_array_out[1][9] .power_up = "low";

dffeas \i_array_out[3][9] (
	.clk(clk),
	.d(\Mux70~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(i_array_out_9_3),
	.prn(vcc));
defparam \i_array_out[3][9] .is_wysiwyg = "true";
defparam \i_array_out[3][9] .power_up = "low";

cycloneive_lcell_comb \Mux22~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_2),
	.datac(ram_in_reg_5_2),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
defparam \Mux22~0 .lut_mask = 16'hFAFC;
defparam \Mux22~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~1 (
	.dataa(ram_in_reg_6_2),
	.datab(ram_in_reg_7_2),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
defparam \Mux20~1 .lut_mask = 16'hAACC;
defparam \Mux20~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux22~1 (
	.dataa(\Mux22~0_combout ),
	.datab(\Mux20~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
defparam \Mux22~1 .lut_mask = 16'hEEFF;
defparam \Mux22~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_0),
	.datac(ram_in_reg_5_0),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFAFC;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(ram_in_reg_6_0),
	.datab(ram_in_reg_7_0),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hAACC;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\Mux2~0_combout ),
	.datab(\Mux0~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hEEFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux23~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_2),
	.datac(ram_in_reg_4_2),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
defparam \Mux23~0 .lut_mask = 16'hFAFC;
defparam \Mux23~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~0 (
	.dataa(ram_in_reg_5_2),
	.datab(ram_in_reg_6_2),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
defparam \Mux20~0 .lut_mask = 16'hAACC;
defparam \Mux20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux23~1 (
	.dataa(\Mux23~0_combout ),
	.datab(\Mux20~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
defparam \Mux23~1 .lut_mask = 16'hEEFF;
defparam \Mux23~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_0),
	.datac(ram_in_reg_4_0),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFAFC;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(ram_in_reg_5_0),
	.datab(ram_in_reg_6_0),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hAACC;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\Mux3~0_combout ),
	.datab(\Mux0~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hEEFF;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux24~0 (
	.dataa(ram_in_reg_3_2),
	.datab(ram_in_reg_5_2),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
defparam \Mux24~0 .lut_mask = 16'hACFF;
defparam \Mux24~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux25~0 (
	.dataa(ram_in_reg_2_2),
	.datab(ram_in_reg_4_2),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
defparam \Mux25~0 .lut_mask = 16'hAACC;
defparam \Mux25~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux24~1 (
	.dataa(\Mux24~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux25~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
defparam \Mux24~1 .lut_mask = 16'hFEFE;
defparam \Mux24~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(ram_in_reg_3_0),
	.datab(ram_in_reg_5_0),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hACFF;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(ram_in_reg_2_0),
	.datab(ram_in_reg_4_0),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hAACC;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\Mux4~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux5~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFEFE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~0 (
	.dataa(ram_in_reg_1_2),
	.datab(ram_in_reg_3_2),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
defparam \Mux26~0 .lut_mask = 16'hAACC;
defparam \Mux26~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux25~1 (
	.dataa(\Mux26~0_combout ),
	.datab(\Mux25~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
defparam \Mux25~1 .lut_mask = 16'hAACC;
defparam \Mux25~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(ram_in_reg_1_0),
	.datab(ram_in_reg_3_0),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hAACC;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux6~0_combout ),
	.datab(\Mux5~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hAACC;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~1 (
	.dataa(ram_in_reg_0_2),
	.datab(ram_in_reg_2_2),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
defparam \Mux26~1 .lut_mask = 16'hAACC;
defparam \Mux26~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux26~2 (
	.dataa(\Mux26~1_combout ),
	.datab(\Mux26~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
defparam \Mux26~2 .lut_mask = 16'hAACC;
defparam \Mux26~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(ram_in_reg_0_0),
	.datab(ram_in_reg_2_0),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hAACC;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(\Mux6~1_combout ),
	.datab(\Mux6~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hAACC;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux27~0 (
	.dataa(\Mux26~1_combout ),
	.datab(ram_in_reg_1_2),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
defparam \Mux27~0 .lut_mask = 16'hACFF;
defparam \Mux27~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(\Mux6~1_combout ),
	.datab(ram_in_reg_1_0),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hACFF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux32~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_3),
	.datac(ram_in_reg_5_3),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
defparam \Mux32~0 .lut_mask = 16'hFAFC;
defparam \Mux32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~1 (
	.dataa(ram_in_reg_6_3),
	.datab(ram_in_reg_7_3),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
defparam \Mux30~1 .lut_mask = 16'hAACC;
defparam \Mux30~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux32~1 (
	.dataa(\Mux32~0_combout ),
	.datab(\Mux30~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
defparam \Mux32~1 .lut_mask = 16'hEEFF;
defparam \Mux32~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_1),
	.datac(ram_in_reg_5_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFAFC;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~1 (
	.dataa(ram_in_reg_6_1),
	.datab(ram_in_reg_7_1),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
defparam \Mux10~1 .lut_mask = 16'hAACC;
defparam \Mux10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~1 (
	.dataa(\Mux12~0_combout ),
	.datab(\Mux10~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
defparam \Mux12~1 .lut_mask = 16'hEEFF;
defparam \Mux12~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux33~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_3),
	.datac(ram_in_reg_4_3),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
defparam \Mux33~0 .lut_mask = 16'hFAFC;
defparam \Mux33~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(ram_in_reg_5_3),
	.datab(ram_in_reg_6_3),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hAACC;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux33~1 (
	.dataa(\Mux33~0_combout ),
	.datab(\Mux30~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
defparam \Mux33~1 .lut_mask = 16'hEEFF;
defparam \Mux33~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_1),
	.datac(ram_in_reg_4_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFAFC;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~0 (
	.dataa(ram_in_reg_5_1),
	.datab(ram_in_reg_6_1),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hAACC;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~1 (
	.dataa(\Mux13~0_combout ),
	.datab(\Mux10~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
defparam \Mux13~1 .lut_mask = 16'hEEFF;
defparam \Mux13~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux34~0 (
	.dataa(ram_in_reg_3_3),
	.datab(ram_in_reg_5_3),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
defparam \Mux34~0 .lut_mask = 16'hACFF;
defparam \Mux34~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux35~0 (
	.dataa(ram_in_reg_2_3),
	.datab(ram_in_reg_4_3),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
defparam \Mux35~0 .lut_mask = 16'hAACC;
defparam \Mux35~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux34~1 (
	.dataa(\Mux34~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux35~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
defparam \Mux34~1 .lut_mask = 16'hFEFE;
defparam \Mux34~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~0 (
	.dataa(ram_in_reg_3_1),
	.datab(ram_in_reg_5_1),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
defparam \Mux14~0 .lut_mask = 16'hACFF;
defparam \Mux14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(ram_in_reg_2_1),
	.datab(ram_in_reg_4_1),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAACC;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~1 (
	.dataa(\Mux14~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux15~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
defparam \Mux14~1 .lut_mask = 16'hFEFE;
defparam \Mux14~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux36~0 (
	.dataa(ram_in_reg_1_3),
	.datab(ram_in_reg_3_3),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
defparam \Mux36~0 .lut_mask = 16'hAACC;
defparam \Mux36~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux35~1 (
	.dataa(\Mux36~0_combout ),
	.datab(\Mux35~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
defparam \Mux35~1 .lut_mask = 16'hAACC;
defparam \Mux35~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(ram_in_reg_1_1),
	.datab(ram_in_reg_3_1),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hAACC;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~1 (
	.dataa(\Mux16~0_combout ),
	.datab(\Mux15~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
defparam \Mux15~1 .lut_mask = 16'hAACC;
defparam \Mux15~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux36~1 (
	.dataa(ram_in_reg_0_3),
	.datab(ram_in_reg_2_3),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
defparam \Mux36~1 .lut_mask = 16'hAACC;
defparam \Mux36~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux36~2 (
	.dataa(\Mux36~1_combout ),
	.datab(\Mux36~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
defparam \Mux36~2 .lut_mask = 16'hAACC;
defparam \Mux36~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~1 (
	.dataa(ram_in_reg_0_1),
	.datab(ram_in_reg_2_1),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hAACC;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~2 (
	.dataa(\Mux16~1_combout ),
	.datab(\Mux16~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
defparam \Mux16~2 .lut_mask = 16'hAACC;
defparam \Mux16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux37~0 (
	.dataa(\Mux36~1_combout ),
	.datab(ram_in_reg_1_3),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'hACFF;
defparam \Mux37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux17~0 (
	.dataa(\Mux16~1_combout ),
	.datab(ram_in_reg_1_1),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'hACFF;
defparam \Mux17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux62~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_6),
	.datac(ram_in_reg_5_6),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
defparam \Mux62~0 .lut_mask = 16'hFAFC;
defparam \Mux62~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux60~1 (
	.dataa(ram_in_reg_6_6),
	.datab(ram_in_reg_7_6),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
defparam \Mux60~1 .lut_mask = 16'hAACC;
defparam \Mux60~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux62~1 (
	.dataa(\Mux62~0_combout ),
	.datab(\Mux60~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
defparam \Mux62~1 .lut_mask = 16'hEEFF;
defparam \Mux62~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux42~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_4),
	.datac(ram_in_reg_5_4),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
defparam \Mux42~0 .lut_mask = 16'hFAFC;
defparam \Mux42~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux40~1 (
	.dataa(ram_in_reg_6_4),
	.datab(ram_in_reg_7_4),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
defparam \Mux40~1 .lut_mask = 16'hAACC;
defparam \Mux40~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux42~1 (
	.dataa(\Mux42~0_combout ),
	.datab(\Mux40~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
defparam \Mux42~1 .lut_mask = 16'hEEFF;
defparam \Mux42~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux63~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_6),
	.datac(ram_in_reg_4_6),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
defparam \Mux63~0 .lut_mask = 16'hFAFC;
defparam \Mux63~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux60~0 (
	.dataa(ram_in_reg_5_6),
	.datab(ram_in_reg_6_6),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
defparam \Mux60~0 .lut_mask = 16'hAACC;
defparam \Mux60~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux63~1 (
	.dataa(\Mux63~0_combout ),
	.datab(\Mux60~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
defparam \Mux63~1 .lut_mask = 16'hEEFF;
defparam \Mux63~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux43~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_4),
	.datac(ram_in_reg_4_4),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
defparam \Mux43~0 .lut_mask = 16'hFAFC;
defparam \Mux43~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux40~0 (
	.dataa(ram_in_reg_5_4),
	.datab(ram_in_reg_6_4),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
defparam \Mux40~0 .lut_mask = 16'hAACC;
defparam \Mux40~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux43~1 (
	.dataa(\Mux43~0_combout ),
	.datab(\Mux40~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
defparam \Mux43~1 .lut_mask = 16'hEEFF;
defparam \Mux43~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux64~0 (
	.dataa(ram_in_reg_3_6),
	.datab(ram_in_reg_5_6),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux64~0_combout ),
	.cout());
defparam \Mux64~0 .lut_mask = 16'hACFF;
defparam \Mux64~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux65~0 (
	.dataa(ram_in_reg_2_6),
	.datab(ram_in_reg_4_6),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux65~0_combout ),
	.cout());
defparam \Mux65~0 .lut_mask = 16'hAACC;
defparam \Mux65~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux64~1 (
	.dataa(\Mux64~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux65~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux64~1_combout ),
	.cout());
defparam \Mux64~1 .lut_mask = 16'hFEFE;
defparam \Mux64~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux44~0 (
	.dataa(ram_in_reg_3_4),
	.datab(ram_in_reg_5_4),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
defparam \Mux44~0 .lut_mask = 16'hACFF;
defparam \Mux44~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux45~0 (
	.dataa(ram_in_reg_2_4),
	.datab(ram_in_reg_4_4),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
defparam \Mux45~0 .lut_mask = 16'hAACC;
defparam \Mux45~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux44~1 (
	.dataa(\Mux44~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux45~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
defparam \Mux44~1 .lut_mask = 16'hFEFE;
defparam \Mux44~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux66~0 (
	.dataa(ram_in_reg_1_6),
	.datab(ram_in_reg_3_6),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux66~0_combout ),
	.cout());
defparam \Mux66~0 .lut_mask = 16'hAACC;
defparam \Mux66~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux65~1 (
	.dataa(\Mux66~0_combout ),
	.datab(\Mux65~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux65~1_combout ),
	.cout());
defparam \Mux65~1 .lut_mask = 16'hAACC;
defparam \Mux65~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux46~0 (
	.dataa(ram_in_reg_1_4),
	.datab(ram_in_reg_3_4),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
defparam \Mux46~0 .lut_mask = 16'hAACC;
defparam \Mux46~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux45~1 (
	.dataa(\Mux46~0_combout ),
	.datab(\Mux45~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
defparam \Mux45~1 .lut_mask = 16'hAACC;
defparam \Mux45~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux66~1 (
	.dataa(ram_in_reg_0_6),
	.datab(ram_in_reg_2_6),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux66~1_combout ),
	.cout());
defparam \Mux66~1 .lut_mask = 16'hAACC;
defparam \Mux66~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux66~2 (
	.dataa(\Mux66~1_combout ),
	.datab(\Mux66~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux66~2_combout ),
	.cout());
defparam \Mux66~2 .lut_mask = 16'hAACC;
defparam \Mux66~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux46~1 (
	.dataa(ram_in_reg_0_4),
	.datab(ram_in_reg_2_4),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
defparam \Mux46~1 .lut_mask = 16'hAACC;
defparam \Mux46~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux46~2 (
	.dataa(\Mux46~1_combout ),
	.datab(\Mux46~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
defparam \Mux46~2 .lut_mask = 16'hAACC;
defparam \Mux46~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux67~0 (
	.dataa(\Mux66~1_combout ),
	.datab(ram_in_reg_1_6),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux67~0_combout ),
	.cout());
defparam \Mux67~0 .lut_mask = 16'hACFF;
defparam \Mux67~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux47~0 (
	.dataa(\Mux46~1_combout ),
	.datab(ram_in_reg_1_4),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
defparam \Mux47~0 .lut_mask = 16'hACFF;
defparam \Mux47~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux72~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_7),
	.datac(ram_in_reg_5_7),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux72~0_combout ),
	.cout());
defparam \Mux72~0 .lut_mask = 16'hFAFC;
defparam \Mux72~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux70~1 (
	.dataa(ram_in_reg_6_7),
	.datab(ram_in_reg_7_7),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux70~1_combout ),
	.cout());
defparam \Mux70~1 .lut_mask = 16'hAACC;
defparam \Mux70~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux72~1 (
	.dataa(\Mux72~0_combout ),
	.datab(\Mux70~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux72~1_combout ),
	.cout());
defparam \Mux72~1 .lut_mask = 16'hEEFF;
defparam \Mux72~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux52~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_4_5),
	.datac(ram_in_reg_5_5),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
defparam \Mux52~0 .lut_mask = 16'hFAFC;
defparam \Mux52~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux50~1 (
	.dataa(ram_in_reg_6_5),
	.datab(ram_in_reg_7_5),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
defparam \Mux50~1 .lut_mask = 16'hAACC;
defparam \Mux50~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux52~1 (
	.dataa(\Mux52~0_combout ),
	.datab(\Mux50~1_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
defparam \Mux52~1 .lut_mask = 16'hEEFF;
defparam \Mux52~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux73~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_7),
	.datac(ram_in_reg_4_7),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux73~0_combout ),
	.cout());
defparam \Mux73~0 .lut_mask = 16'hFAFC;
defparam \Mux73~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux70~0 (
	.dataa(ram_in_reg_5_7),
	.datab(ram_in_reg_6_7),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux70~0_combout ),
	.cout());
defparam \Mux70~0 .lut_mask = 16'hAACC;
defparam \Mux70~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux73~1 (
	.dataa(\Mux73~0_combout ),
	.datab(\Mux70~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux73~1_combout ),
	.cout());
defparam \Mux73~1 .lut_mask = 16'hEEFF;
defparam \Mux73~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux53~0 (
	.dataa(slb_last_1),
	.datab(ram_in_reg_3_5),
	.datac(ram_in_reg_4_5),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
defparam \Mux53~0 .lut_mask = 16'hFAFC;
defparam \Mux53~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux50~0 (
	.dataa(ram_in_reg_5_5),
	.datab(ram_in_reg_6_5),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
defparam \Mux50~0 .lut_mask = 16'hAACC;
defparam \Mux50~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux53~1 (
	.dataa(\Mux53~0_combout ),
	.datab(\Mux50~0_combout ),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
defparam \Mux53~1 .lut_mask = 16'hEEFF;
defparam \Mux53~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux74~0 (
	.dataa(ram_in_reg_3_7),
	.datab(ram_in_reg_5_7),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux74~0_combout ),
	.cout());
defparam \Mux74~0 .lut_mask = 16'hACFF;
defparam \Mux74~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux75~0 (
	.dataa(ram_in_reg_2_7),
	.datab(ram_in_reg_4_7),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux75~0_combout ),
	.cout());
defparam \Mux75~0 .lut_mask = 16'hAACC;
defparam \Mux75~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux74~1 (
	.dataa(\Mux74~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux75~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux74~1_combout ),
	.cout());
defparam \Mux74~1 .lut_mask = 16'hFEFE;
defparam \Mux74~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux54~0 (
	.dataa(ram_in_reg_3_5),
	.datab(ram_in_reg_5_5),
	.datac(slb_last_1),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
defparam \Mux54~0 .lut_mask = 16'hACFF;
defparam \Mux54~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux55~0 (
	.dataa(ram_in_reg_2_5),
	.datab(ram_in_reg_4_5),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
defparam \Mux55~0 .lut_mask = 16'hAACC;
defparam \Mux55~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux54~1 (
	.dataa(\Mux54~0_combout ),
	.datab(slb_last_0),
	.datac(\Mux55~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
defparam \Mux54~1 .lut_mask = 16'hFEFE;
defparam \Mux54~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux76~0 (
	.dataa(ram_in_reg_1_7),
	.datab(ram_in_reg_3_7),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux76~0_combout ),
	.cout());
defparam \Mux76~0 .lut_mask = 16'hAACC;
defparam \Mux76~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux75~1 (
	.dataa(\Mux76~0_combout ),
	.datab(\Mux75~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux75~1_combout ),
	.cout());
defparam \Mux75~1 .lut_mask = 16'hAACC;
defparam \Mux75~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux56~0 (
	.dataa(ram_in_reg_1_5),
	.datab(ram_in_reg_3_5),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
defparam \Mux56~0 .lut_mask = 16'hAACC;
defparam \Mux56~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux55~1 (
	.dataa(\Mux56~0_combout ),
	.datab(\Mux55~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
defparam \Mux55~1 .lut_mask = 16'hAACC;
defparam \Mux55~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux76~1 (
	.dataa(ram_in_reg_0_7),
	.datab(ram_in_reg_2_7),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux76~1_combout ),
	.cout());
defparam \Mux76~1 .lut_mask = 16'hAACC;
defparam \Mux76~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux76~2 (
	.dataa(\Mux76~1_combout ),
	.datab(\Mux76~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux76~2_combout ),
	.cout());
defparam \Mux76~2 .lut_mask = 16'hAACC;
defparam \Mux76~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux56~1 (
	.dataa(ram_in_reg_0_5),
	.datab(ram_in_reg_2_5),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
defparam \Mux56~1 .lut_mask = 16'hAACC;
defparam \Mux56~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux56~2 (
	.dataa(\Mux56~1_combout ),
	.datab(\Mux56~0_combout ),
	.datac(gnd),
	.datad(slb_last_0),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
defparam \Mux56~2 .lut_mask = 16'hAACC;
defparam \Mux56~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux77~0 (
	.dataa(\Mux76~1_combout ),
	.datab(ram_in_reg_1_7),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux77~0_combout ),
	.cout());
defparam \Mux77~0 .lut_mask = 16'hACFF;
defparam \Mux77~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux57~0 (
	.dataa(\Mux56~1_combout ),
	.datab(ram_in_reg_1_5),
	.datac(slb_last_0),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
defparam \Mux57~0 .lut_mask = 16'hACFF;
defparam \Mux57~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_array_out[2][9]~0 (
	.dataa(slb_last_2),
	.datab(slb_last_0),
	.datac(gnd),
	.datad(slb_last_1),
	.cin(gnd),
	.combout(\i_array_out[2][9]~0_combout ),
	.cout());
defparam \i_array_out[2][9]~0 .lut_mask = 16'hEEFF;
defparam \i_array_out[2][9]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_array_out[2][9]~1 (
	.dataa(slb_last_1),
	.datab(slb_last_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\i_array_out[2][9]~1_combout ),
	.cout());
defparam \i_array_out[2][9]~1 .lut_mask = 16'hEEEE;
defparam \i_array_out[2][9]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_8_0),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(ram_in_reg_7_0),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux1~0_combout ),
	.datad(ram_in_reg_4_0),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux21~0 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux20~0_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_8_2),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
defparam \Mux21~0 .lut_mask = 16'hFFDE;
defparam \Mux21~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux21~1 (
	.dataa(ram_in_reg_7_2),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux21~0_combout ),
	.datad(ram_in_reg_4_2),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
defparam \Mux21~1 .lut_mask = 16'hFFBE;
defparam \Mux21~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~0 (
	.dataa(ram_in_reg_0_0),
	.datab(ram_in_reg_1_0),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hACFF;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux28~0 (
	.dataa(ram_in_reg_0_2),
	.datab(ram_in_reg_1_2),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
defparam \Mux28~0 .lut_mask = 16'hACFF;
defparam \Mux28~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(ram_in_reg_0_0),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hBFFF;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux29~0 (
	.dataa(ram_in_reg_0_2),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
defparam \Mux29~0 .lut_mask = 16'hBFFF;
defparam \Mux29~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux10~0_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_8_1),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hFFDE;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~1 (
	.dataa(ram_in_reg_7_1),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux11~0_combout ),
	.datad(ram_in_reg_4_1),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
defparam \Mux11~1 .lut_mask = 16'hFFBE;
defparam \Mux11~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux31~0 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux30~0_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_8_3),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hFFDE;
defparam \Mux31~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux31~1 (
	.dataa(ram_in_reg_7_3),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux31~0_combout ),
	.datad(ram_in_reg_4_3),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
defparam \Mux31~1 .lut_mask = 16'hFFBE;
defparam \Mux31~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux18~0 (
	.dataa(ram_in_reg_0_1),
	.datab(ram_in_reg_1_1),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
defparam \Mux18~0 .lut_mask = 16'hACFF;
defparam \Mux18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux38~0 (
	.dataa(ram_in_reg_0_3),
	.datab(ram_in_reg_1_3),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
defparam \Mux38~0 .lut_mask = 16'hACFF;
defparam \Mux38~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux19~0 (
	.dataa(ram_in_reg_0_1),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
defparam \Mux19~0 .lut_mask = 16'hBFFF;
defparam \Mux19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux39~0 (
	.dataa(ram_in_reg_0_3),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
defparam \Mux39~0 .lut_mask = 16'hBFFF;
defparam \Mux39~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux0~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_0),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFDE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(ram_in_reg_8_0),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux0~2_combout ),
	.datad(ram_in_reg_5_0),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFBE;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux20~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_2),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
defparam \Mux20~2 .lut_mask = 16'hFFDE;
defparam \Mux20~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux20~3 (
	.dataa(ram_in_reg_8_2),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux20~2_combout ),
	.datad(ram_in_reg_5_2),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
defparam \Mux20~3 .lut_mask = 16'hFFBE;
defparam \Mux20~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux10~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_1),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
defparam \Mux10~2 .lut_mask = 16'hFFDE;
defparam \Mux10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~3 (
	.dataa(ram_in_reg_8_1),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux10~2_combout ),
	.datad(ram_in_reg_5_1),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
defparam \Mux10~3 .lut_mask = 16'hFFBE;
defparam \Mux10~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux30~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_3),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
defparam \Mux30~2 .lut_mask = 16'hFFDE;
defparam \Mux30~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~3 (
	.dataa(ram_in_reg_8_3),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux30~2_combout ),
	.datad(ram_in_reg_5_3),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
defparam \Mux30~3 .lut_mask = 16'hFFBE;
defparam \Mux30~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux41~0 (
	.dataa(\i_array_out[2][9]~1_combout ),
	.datab(ram_in_reg_7_4),
	.datac(\i_array_out[2][9]~0_combout ),
	.datad(ram_in_reg_8_4),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
defparam \Mux41~0 .lut_mask = 16'hFFDE;
defparam \Mux41~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux41~1 (
	.dataa(\Mux40~0_combout ),
	.datab(\i_array_out[2][9]~1_combout ),
	.datac(\Mux41~0_combout ),
	.datad(ram_in_reg_4_4),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
defparam \Mux41~1 .lut_mask = 16'hFFBE;
defparam \Mux41~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux61~0 (
	.dataa(\i_array_out[2][9]~1_combout ),
	.datab(ram_in_reg_7_6),
	.datac(\i_array_out[2][9]~0_combout ),
	.datad(ram_in_reg_8_6),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
defparam \Mux61~0 .lut_mask = 16'hFFDE;
defparam \Mux61~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux61~1 (
	.dataa(\Mux60~0_combout ),
	.datab(\i_array_out[2][9]~1_combout ),
	.datac(\Mux61~0_combout ),
	.datad(ram_in_reg_4_6),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
defparam \Mux61~1 .lut_mask = 16'hFFBE;
defparam \Mux61~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux48~0 (
	.dataa(ram_in_reg_0_4),
	.datab(ram_in_reg_1_4),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
defparam \Mux48~0 .lut_mask = 16'hACFF;
defparam \Mux48~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux68~0 (
	.dataa(ram_in_reg_0_6),
	.datab(ram_in_reg_1_6),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux68~0_combout ),
	.cout());
defparam \Mux68~0 .lut_mask = 16'hACFF;
defparam \Mux68~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux49~0 (
	.dataa(ram_in_reg_0_4),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
defparam \Mux49~0 .lut_mask = 16'hBFFF;
defparam \Mux49~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux69~0 (
	.dataa(ram_in_reg_0_6),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux69~0_combout ),
	.cout());
defparam \Mux69~0 .lut_mask = 16'hBFFF;
defparam \Mux69~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux51~0 (
	.dataa(\i_array_out[2][9]~1_combout ),
	.datab(ram_in_reg_7_5),
	.datac(\i_array_out[2][9]~0_combout ),
	.datad(ram_in_reg_8_5),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
defparam \Mux51~0 .lut_mask = 16'hFFDE;
defparam \Mux51~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux51~1 (
	.dataa(\Mux50~0_combout ),
	.datab(\i_array_out[2][9]~1_combout ),
	.datac(\Mux51~0_combout ),
	.datad(ram_in_reg_4_5),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
defparam \Mux51~1 .lut_mask = 16'hFFBE;
defparam \Mux51~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux71~0 (
	.dataa(\i_array_out[2][9]~1_combout ),
	.datab(ram_in_reg_7_7),
	.datac(\i_array_out[2][9]~0_combout ),
	.datad(ram_in_reg_8_7),
	.cin(gnd),
	.combout(\Mux71~0_combout ),
	.cout());
defparam \Mux71~0 .lut_mask = 16'hFFDE;
defparam \Mux71~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux71~1 (
	.dataa(\Mux70~0_combout ),
	.datab(\i_array_out[2][9]~1_combout ),
	.datac(\Mux71~0_combout ),
	.datad(ram_in_reg_4_7),
	.cin(gnd),
	.combout(\Mux71~1_combout ),
	.cout());
defparam \Mux71~1 .lut_mask = 16'hFFBE;
defparam \Mux71~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux58~0 (
	.dataa(ram_in_reg_0_5),
	.datab(ram_in_reg_1_5),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
defparam \Mux58~0 .lut_mask = 16'hACFF;
defparam \Mux58~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux78~0 (
	.dataa(ram_in_reg_0_7),
	.datab(ram_in_reg_1_7),
	.datac(slb_last_0),
	.datad(\i_array_out[2][9]~1_combout ),
	.cin(gnd),
	.combout(\Mux78~0_combout ),
	.cout());
defparam \Mux78~0 .lut_mask = 16'hACFF;
defparam \Mux78~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux59~0 (
	.dataa(ram_in_reg_0_5),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
defparam \Mux59~0 .lut_mask = 16'hBFFF;
defparam \Mux59~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux79~0 (
	.dataa(ram_in_reg_0_7),
	.datab(slb_last_0),
	.datac(slb_last_1),
	.datad(slb_last_2),
	.cin(gnd),
	.combout(\Mux79~0_combout ),
	.cout());
defparam \Mux79~0 .lut_mask = 16'hBFFF;
defparam \Mux79~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux40~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux40~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_4),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
defparam \Mux40~2 .lut_mask = 16'hFFDE;
defparam \Mux40~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux40~3 (
	.dataa(ram_in_reg_8_4),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux40~2_combout ),
	.datad(ram_in_reg_5_4),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
defparam \Mux40~3 .lut_mask = 16'hFFBE;
defparam \Mux40~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux60~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux60~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_6),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
defparam \Mux60~2 .lut_mask = 16'hFFDE;
defparam \Mux60~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux60~3 (
	.dataa(ram_in_reg_8_6),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux60~2_combout ),
	.datad(ram_in_reg_5_6),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
defparam \Mux60~3 .lut_mask = 16'hFFBE;
defparam \Mux60~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux50~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux50~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_5),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
defparam \Mux50~2 .lut_mask = 16'hFFDE;
defparam \Mux50~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux50~3 (
	.dataa(ram_in_reg_8_5),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux50~2_combout ),
	.datad(ram_in_reg_5_5),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
defparam \Mux50~3 .lut_mask = 16'hFFBE;
defparam \Mux50~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux70~2 (
	.dataa(\i_array_out[2][9]~0_combout ),
	.datab(\Mux70~1_combout ),
	.datac(\i_array_out[2][9]~1_combout ),
	.datad(ram_in_reg_9_7),
	.cin(gnd),
	.combout(\Mux70~2_combout ),
	.cout());
defparam \Mux70~2 .lut_mask = 16'hFFDE;
defparam \Mux70~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux70~3 (
	.dataa(ram_in_reg_8_7),
	.datab(\i_array_out[2][9]~0_combout ),
	.datac(\Mux70~2_combout ),
	.datad(ram_in_reg_5_7),
	.cin(gnd),
	.combout(\Mux70~3_combout ),
	.cout());
defparam \Mux70~3 .lut_mask = 16'hFFBE;
defparam \Mux70~3 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_bfp_o (
	global_clock_enable,
	tdl_arr_0,
	sdetdIDLE,
	slb_i_0,
	slb_i_1,
	slb_i_2,
	slb_i_3,
	Mux2,
	Mux1,
	tdl_arr_6,
	reg_no_twiddle605,
	reg_no_twiddle609,
	reg_no_twiddle615,
	reg_no_twiddle619,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_5_12,
	tdl_arr_9_12,
	tdl_arr_5_13,
	tdl_arr_9_13,
	tdl_arr_5_14,
	tdl_arr_9_14,
	tdl_arr_5_15,
	tdl_arr_9_15,
	reg_no_twiddle606,
	reg_no_twiddle616,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	reg_no_twiddle607,
	reg_no_twiddle617,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_7_12,
	tdl_arr_7_13,
	tdl_arr_7_14,
	tdl_arr_7_15,
	reg_no_twiddle608,
	reg_no_twiddle618,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_8_12,
	tdl_arr_8_13,
	tdl_arr_8_14,
	tdl_arr_8_15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	tdl_arr_0;
output 	sdetdIDLE;
output 	slb_i_0;
output 	slb_i_1;
output 	slb_i_2;
output 	slb_i_3;
output 	Mux2;
output 	Mux1;
input 	tdl_arr_6;
input 	reg_no_twiddle605;
input 	reg_no_twiddle609;
input 	reg_no_twiddle615;
input 	reg_no_twiddle619;
input 	tdl_arr_5_1;
input 	tdl_arr_9_1;
input 	tdl_arr_5_11;
input 	tdl_arr_9_11;
input 	tdl_arr_5_12;
input 	tdl_arr_9_12;
input 	tdl_arr_5_13;
input 	tdl_arr_9_13;
input 	tdl_arr_5_14;
input 	tdl_arr_9_14;
input 	tdl_arr_5_15;
input 	tdl_arr_9_15;
input 	reg_no_twiddle606;
input 	reg_no_twiddle616;
input 	tdl_arr_6_1;
input 	tdl_arr_6_11;
input 	tdl_arr_6_12;
input 	tdl_arr_6_13;
input 	tdl_arr_6_14;
input 	tdl_arr_6_15;
input 	reg_no_twiddle607;
input 	reg_no_twiddle617;
input 	tdl_arr_7_1;
input 	tdl_arr_7_11;
input 	tdl_arr_7_12;
input 	tdl_arr_7_13;
input 	tdl_arr_7_14;
input 	tdl_arr_7_15;
input 	reg_no_twiddle608;
input 	reg_no_twiddle618;
input 	tdl_arr_8_1;
input 	tdl_arr_8_11;
input 	tdl_arr_8_12;
input 	tdl_arr_8_13;
input 	tdl_arr_8_14;
input 	tdl_arr_8_15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_blk_float:gen_b:delay_next_blk|tdl_arr[0]~q ;
wire \gain_lut_8pts~0_combout ;
wire \gain_lut_8pts~1_combout ;
wire \gain_lut_8pts~2_combout ;
wire \gain_lut_8pts~3_combout ;
wire \gain_lut_8pts~4_combout ;
wire \Selector1~0_combout ;
wire \sdetd.SLBI~0_combout ;
wire \sdetd.SLBI~q ;
wire \del_np_cnt[0]~5_combout ;
wire \Selector0~0_combout ;
wire \Equal0~0_combout ;
wire \Selector0~1_combout ;
wire \sdetd.BLOCK_READY~q ;
wire \delay_next_pass4~2_combout ;
wire \del_np_cnt[0]~q ;
wire \del_np_cnt[0]~6 ;
wire \del_np_cnt[1]~7_combout ;
wire \del_np_cnt[1]~q ;
wire \del_np_cnt[1]~8 ;
wire \del_np_cnt[2]~9_combout ;
wire \del_np_cnt[2]~q ;
wire \del_np_cnt[2]~10 ;
wire \del_np_cnt[3]~11_combout ;
wire \del_np_cnt[3]~q ;
wire \del_np_cnt[3]~12 ;
wire \del_np_cnt[4]~13_combout ;
wire \del_np_cnt[4]~q ;
wire \Equal1~0_combout ;
wire \Selector2~0_combout ;
wire \sdetd.DISABLE~q ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \sdetd.ENABLE~q ;
wire \sdetd~8_combout ;
wire \sdetd.GBLK~q ;
wire \gain_lut_8pts~5_combout ;
wire \gain_lut_8pts[0]~q ;
wire \Selector6~0_combout ;
wire \gain_lut_blk[0]~q ;
wire \Selector10~0_combout ;
wire \slb_i[3]~0_combout ;
wire \gain_lut_8pts~6_combout ;
wire \gain_lut_8pts~7_combout ;
wire \gain_lut_8pts~8_combout ;
wire \gain_lut_8pts~9_combout ;
wire \gain_lut_8pts~10_combout ;
wire \gain_lut_8pts~11_combout ;
wire \gain_lut_8pts[1]~q ;
wire \Selector5~0_combout ;
wire \gain_lut_blk[1]~q ;
wire \Selector9~0_combout ;
wire \gain_lut_8pts~12_combout ;
wire \gain_lut_8pts~13_combout ;
wire \gain_lut_8pts~14_combout ;
wire \gain_lut_8pts~15_combout ;
wire \gain_lut_8pts~16_combout ;
wire \gain_lut_8pts~17_combout ;
wire \gain_lut_8pts[2]~q ;
wire \Selector4~0_combout ;
wire \gain_lut_blk[2]~q ;
wire \Selector8~0_combout ;
wire \gain_lut_8pts~18_combout ;
wire \gain_lut_8pts~19_combout ;
wire \gain_lut_8pts~20_combout ;
wire \gain_lut_8pts~21_combout ;
wire \gain_lut_8pts~22_combout ;
wire \gain_lut_8pts~23_combout ;
wire \gain_lut_8pts[3]~q ;
wire \Selector3~0_combout ;
wire \gain_lut_blk[3]~q ;
wire \Selector7~0_combout ;


fftsign_asj_fft_tdl_bit_rst_1 \gen_blk_float:gen_b:delay_next_blk (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(tdl_arr_0),
	.tdl_arr_01(\gen_blk_float:gen_b:delay_next_blk|tdl_arr[0]~q ),
	.clk(clk),
	.reset_n(reset_n));

dffeas \sdetd.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sdetdIDLE),
	.prn(vcc));
defparam \sdetd.IDLE .is_wysiwyg = "true";
defparam \sdetd.IDLE .power_up = "low";

dffeas \slb_i[0] (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_0),
	.prn(vcc));
defparam \slb_i[0] .is_wysiwyg = "true";
defparam \slb_i[0] .power_up = "low";

dffeas \slb_i[1] (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_1),
	.prn(vcc));
defparam \slb_i[1] .is_wysiwyg = "true";
defparam \slb_i[1] .power_up = "low";

dffeas \slb_i[2] (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_2),
	.prn(vcc));
defparam \slb_i[2] .is_wysiwyg = "true";
defparam \slb_i[2] .power_up = "low";

dffeas \slb_i[3] (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_i[3]~0_combout ),
	.q(slb_i_3),
	.prn(vcc));
defparam \slb_i[3] .is_wysiwyg = "true";
defparam \slb_i[3] .power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(slb_i_0),
	.datab(slb_i_1),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(Mux2),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFBFF;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(slb_i_0),
	.datab(slb_i_1),
	.datac(slb_i_2),
	.datad(slb_i_3),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFF;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~0 (
	.dataa(reg_no_twiddle605),
	.datab(reg_no_twiddle609),
	.datac(reg_no_twiddle615),
	.datad(reg_no_twiddle619),
	.cin(gnd),
	.combout(\gain_lut_8pts~0_combout ),
	.cout());
defparam \gain_lut_8pts~0 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~1 (
	.dataa(tdl_arr_5_1),
	.datab(tdl_arr_9_1),
	.datac(tdl_arr_5_11),
	.datad(tdl_arr_9_11),
	.cin(gnd),
	.combout(\gain_lut_8pts~1_combout ),
	.cout());
defparam \gain_lut_8pts~1 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~2 (
	.dataa(tdl_arr_5_12),
	.datab(tdl_arr_9_12),
	.datac(tdl_arr_5_13),
	.datad(tdl_arr_9_13),
	.cin(gnd),
	.combout(\gain_lut_8pts~2_combout ),
	.cout());
defparam \gain_lut_8pts~2 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~3 (
	.dataa(tdl_arr_5_14),
	.datab(tdl_arr_9_14),
	.datac(tdl_arr_5_15),
	.datad(tdl_arr_9_15),
	.cin(gnd),
	.combout(\gain_lut_8pts~3_combout ),
	.cout());
defparam \gain_lut_8pts~3 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~4 (
	.dataa(\gain_lut_8pts~0_combout ),
	.datab(\gain_lut_8pts~1_combout ),
	.datac(\gain_lut_8pts~2_combout ),
	.datad(\gain_lut_8pts~3_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~4_combout ),
	.cout());
defparam \gain_lut_8pts~4 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\sdetd.ENABLE~q ),
	.datab(tdl_arr_6),
	.datac(\gen_blk_float:gen_b:delay_next_blk|tdl_arr[0]~q ),
	.datad(sdetdIDLE),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hBFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sdetd.SLBI~0 (
	.dataa(reset_n),
	.datab(\sdetd.GBLK~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sdetd.SLBI~0_combout ),
	.cout());
defparam \sdetd.SLBI~0 .lut_mask = 16'hEEEE;
defparam \sdetd.SLBI~0 .sum_lutc_input = "datac";

dffeas \sdetd.SLBI (
	.clk(clk),
	.d(\sdetd.SLBI~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdetd.SLBI~q ),
	.prn(vcc));
defparam \sdetd.SLBI .is_wysiwyg = "true";
defparam \sdetd.SLBI .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[0]~5 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_np_cnt[0]~5_combout ),
	.cout(\del_np_cnt[0]~6 ));
defparam \del_np_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \del_np_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\sdetd.ENABLE~q ),
	.datab(\gen_blk_float:gen_b:delay_next_blk|tdl_arr[0]~q ),
	.datac(gnd),
	.datad(tdl_arr_6),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEEFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(\del_np_cnt[2]~q ),
	.datac(\del_np_cnt[1]~q ),
	.datad(\del_np_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(\Selector0~0_combout ),
	.datab(\sdetd.BLOCK_READY~q ),
	.datac(\del_np_cnt[4]~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hEFFF;
defparam \Selector0~1 .sum_lutc_input = "datac";

dffeas \sdetd.BLOCK_READY (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdetd.BLOCK_READY~q ),
	.prn(vcc));
defparam \sdetd.BLOCK_READY .is_wysiwyg = "true";
defparam \sdetd.BLOCK_READY .power_up = "low";

cycloneive_lcell_comb \delay_next_pass4~2 (
	.dataa(\sdetd.DISABLE~q ),
	.datab(\sdetd.BLOCK_READY~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\delay_next_pass4~2_combout ),
	.cout());
defparam \delay_next_pass4~2 .lut_mask = 16'h7777;
defparam \delay_next_pass4~2 .sum_lutc_input = "datac";

dffeas \del_np_cnt[0] (
	.clk(clk),
	.d(\del_np_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass4~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[0]~q ),
	.prn(vcc));
defparam \del_np_cnt[0] .is_wysiwyg = "true";
defparam \del_np_cnt[0] .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[1]~7 (
	.dataa(\del_np_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[0]~6 ),
	.combout(\del_np_cnt[1]~7_combout ),
	.cout(\del_np_cnt[1]~8 ));
defparam \del_np_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[1]~7 .sum_lutc_input = "cin";

dffeas \del_np_cnt[1] (
	.clk(clk),
	.d(\del_np_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass4~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[1]~q ),
	.prn(vcc));
defparam \del_np_cnt[1] .is_wysiwyg = "true";
defparam \del_np_cnt[1] .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[2]~9 (
	.dataa(\del_np_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[1]~8 ),
	.combout(\del_np_cnt[2]~9_combout ),
	.cout(\del_np_cnt[2]~10 ));
defparam \del_np_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \del_np_cnt[2]~9 .sum_lutc_input = "cin";

dffeas \del_np_cnt[2] (
	.clk(clk),
	.d(\del_np_cnt[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass4~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[2]~q ),
	.prn(vcc));
defparam \del_np_cnt[2] .is_wysiwyg = "true";
defparam \del_np_cnt[2] .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[3]~11 (
	.dataa(\del_np_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_np_cnt[2]~10 ),
	.combout(\del_np_cnt[3]~11_combout ),
	.cout(\del_np_cnt[3]~12 ));
defparam \del_np_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \del_np_cnt[3]~11 .sum_lutc_input = "cin";

dffeas \del_np_cnt[3] (
	.clk(clk),
	.d(\del_np_cnt[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass4~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[3]~q ),
	.prn(vcc));
defparam \del_np_cnt[3] .is_wysiwyg = "true";
defparam \del_np_cnt[3] .power_up = "low";

cycloneive_lcell_comb \del_np_cnt[4]~13 (
	.dataa(\del_np_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_np_cnt[3]~12 ),
	.combout(\del_np_cnt[4]~13_combout ),
	.cout());
defparam \del_np_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \del_np_cnt[4]~13 .sum_lutc_input = "cin";

dffeas \del_np_cnt[4] (
	.clk(clk),
	.d(\del_np_cnt[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\delay_next_pass4~2_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_np_cnt[4]~q ),
	.prn(vcc));
defparam \del_np_cnt[4] .is_wysiwyg = "true";
defparam \del_np_cnt[4] .power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\del_np_cnt[0]~q ),
	.datab(\del_np_cnt[1]~q ),
	.datac(\del_np_cnt[3]~q ),
	.datad(\del_np_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\sdetd.SLBI~q ),
	.datab(\sdetd.DISABLE~q ),
	.datac(\del_np_cnt[4]~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \sdetd.DISABLE (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdetd.DISABLE~q ),
	.prn(vcc));
defparam \sdetd.DISABLE .is_wysiwyg = "true";
defparam \sdetd.DISABLE .power_up = "low";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\Selector1~0_combout ),
	.datab(\sdetd.DISABLE~q ),
	.datac(\Equal1~0_combout ),
	.datad(\del_np_cnt[4]~q ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hFEFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\Selector1~1_combout ),
	.datab(\del_np_cnt[4]~q ),
	.datac(\sdetd.BLOCK_READY~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hFFFE;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \sdetd.ENABLE (
	.clk(clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdetd.ENABLE~q ),
	.prn(vcc));
defparam \sdetd.ENABLE .is_wysiwyg = "true";
defparam \sdetd.ENABLE .power_up = "low";

cycloneive_lcell_comb \sdetd~8 (
	.dataa(reset_n),
	.datab(\sdetd.ENABLE~q ),
	.datac(tdl_arr_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\sdetd~8_combout ),
	.cout());
defparam \sdetd~8 .lut_mask = 16'hFEFE;
defparam \sdetd~8 .sum_lutc_input = "datac";

dffeas \sdetd.GBLK (
	.clk(clk),
	.d(\sdetd~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sdetd.GBLK~q ),
	.prn(vcc));
defparam \sdetd.GBLK .is_wysiwyg = "true";
defparam \sdetd.GBLK .power_up = "low";

cycloneive_lcell_comb \gain_lut_8pts~5 (
	.dataa(\gain_lut_8pts~4_combout ),
	.datab(\sdetd.GBLK~q ),
	.datac(\sdetd.ENABLE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~5_combout ),
	.cout());
defparam \gain_lut_8pts~5 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~5 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[0] (
	.clk(clk),
	.d(\gain_lut_8pts~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[0]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[0] .is_wysiwyg = "true";
defparam \gain_lut_8pts[0] .power_up = "low";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\gain_lut_8pts[0]~q ),
	.datab(\gain_lut_blk[0]~q ),
	.datac(\sdetd.GBLK~q ),
	.datad(\sdetd.ENABLE~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hFFFE;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[0] (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[0]~q ),
	.prn(vcc));
defparam \gain_lut_blk[0] .is_wysiwyg = "true";
defparam \gain_lut_blk[0] .power_up = "low";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(\gain_lut_8pts[0]~q ),
	.datab(\gain_lut_blk[0]~q ),
	.datac(gnd),
	.datad(\sdetd.SLBI~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hEEFF;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \slb_i[3]~0 (
	.dataa(global_clock_enable),
	.datab(\sdetd.DISABLE~q ),
	.datac(\sdetd.GBLK~q ),
	.datad(\sdetd.ENABLE~q ),
	.cin(gnd),
	.combout(\slb_i[3]~0_combout ),
	.cout());
defparam \slb_i[3]~0 .lut_mask = 16'hBFFF;
defparam \slb_i[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~6 (
	.dataa(reg_no_twiddle609),
	.datab(reg_no_twiddle606),
	.datac(reg_no_twiddle619),
	.datad(reg_no_twiddle616),
	.cin(gnd),
	.combout(\gain_lut_8pts~6_combout ),
	.cout());
defparam \gain_lut_8pts~6 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~7 (
	.dataa(tdl_arr_9_1),
	.datab(tdl_arr_6_1),
	.datac(tdl_arr_9_11),
	.datad(tdl_arr_6_11),
	.cin(gnd),
	.combout(\gain_lut_8pts~7_combout ),
	.cout());
defparam \gain_lut_8pts~7 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~8 (
	.dataa(tdl_arr_9_12),
	.datab(tdl_arr_6_12),
	.datac(tdl_arr_9_13),
	.datad(tdl_arr_6_13),
	.cin(gnd),
	.combout(\gain_lut_8pts~8_combout ),
	.cout());
defparam \gain_lut_8pts~8 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~9 (
	.dataa(tdl_arr_9_14),
	.datab(tdl_arr_6_14),
	.datac(tdl_arr_9_15),
	.datad(tdl_arr_6_15),
	.cin(gnd),
	.combout(\gain_lut_8pts~9_combout ),
	.cout());
defparam \gain_lut_8pts~9 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~10 (
	.dataa(\gain_lut_8pts~6_combout ),
	.datab(\gain_lut_8pts~7_combout ),
	.datac(\gain_lut_8pts~8_combout ),
	.datad(\gain_lut_8pts~9_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~10_combout ),
	.cout());
defparam \gain_lut_8pts~10 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~11 (
	.dataa(\gain_lut_8pts~10_combout ),
	.datab(\sdetd.GBLK~q ),
	.datac(\sdetd.ENABLE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~11_combout ),
	.cout());
defparam \gain_lut_8pts~11 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~11 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[1] (
	.clk(clk),
	.d(\gain_lut_8pts~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[1]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[1] .is_wysiwyg = "true";
defparam \gain_lut_8pts[1] .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\sdetd.GBLK~q ),
	.datab(\sdetd.ENABLE~q ),
	.datac(\gain_lut_8pts[1]~q ),
	.datad(\gain_lut_blk[1]~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hFFFE;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[1] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[1]~q ),
	.prn(vcc));
defparam \gain_lut_blk[1] .is_wysiwyg = "true";
defparam \gain_lut_blk[1] .power_up = "low";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(\gain_lut_8pts[1]~q ),
	.datab(\gain_lut_blk[1]~q ),
	.datac(gnd),
	.datad(\sdetd.SLBI~q ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hEEFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~12 (
	.dataa(reg_no_twiddle609),
	.datab(reg_no_twiddle607),
	.datac(reg_no_twiddle619),
	.datad(reg_no_twiddle617),
	.cin(gnd),
	.combout(\gain_lut_8pts~12_combout ),
	.cout());
defparam \gain_lut_8pts~12 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~13 (
	.dataa(tdl_arr_9_1),
	.datab(tdl_arr_7_1),
	.datac(tdl_arr_9_11),
	.datad(tdl_arr_7_11),
	.cin(gnd),
	.combout(\gain_lut_8pts~13_combout ),
	.cout());
defparam \gain_lut_8pts~13 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~14 (
	.dataa(tdl_arr_9_12),
	.datab(tdl_arr_7_12),
	.datac(tdl_arr_9_13),
	.datad(tdl_arr_7_13),
	.cin(gnd),
	.combout(\gain_lut_8pts~14_combout ),
	.cout());
defparam \gain_lut_8pts~14 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~15 (
	.dataa(tdl_arr_9_14),
	.datab(tdl_arr_7_14),
	.datac(tdl_arr_9_15),
	.datad(tdl_arr_7_15),
	.cin(gnd),
	.combout(\gain_lut_8pts~15_combout ),
	.cout());
defparam \gain_lut_8pts~15 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~16 (
	.dataa(\gain_lut_8pts~12_combout ),
	.datab(\gain_lut_8pts~13_combout ),
	.datac(\gain_lut_8pts~14_combout ),
	.datad(\gain_lut_8pts~15_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~16_combout ),
	.cout());
defparam \gain_lut_8pts~16 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~17 (
	.dataa(\gain_lut_8pts~16_combout ),
	.datab(\sdetd.GBLK~q ),
	.datac(\sdetd.ENABLE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~17_combout ),
	.cout());
defparam \gain_lut_8pts~17 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~17 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[2] (
	.clk(clk),
	.d(\gain_lut_8pts~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[2]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[2] .is_wysiwyg = "true";
defparam \gain_lut_8pts[2] .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\sdetd.GBLK~q ),
	.datab(\sdetd.ENABLE~q ),
	.datac(\gain_lut_8pts[2]~q ),
	.datad(\gain_lut_blk[2]~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFFFE;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[2] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[2]~q ),
	.prn(vcc));
defparam \gain_lut_blk[2] .is_wysiwyg = "true";
defparam \gain_lut_blk[2] .power_up = "low";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\gain_lut_8pts[2]~q ),
	.datab(\gain_lut_blk[2]~q ),
	.datac(gnd),
	.datad(\sdetd.SLBI~q ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hEEFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~18 (
	.dataa(reg_no_twiddle609),
	.datab(reg_no_twiddle608),
	.datac(reg_no_twiddle619),
	.datad(reg_no_twiddle618),
	.cin(gnd),
	.combout(\gain_lut_8pts~18_combout ),
	.cout());
defparam \gain_lut_8pts~18 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~19 (
	.dataa(tdl_arr_9_1),
	.datab(tdl_arr_8_1),
	.datac(tdl_arr_9_11),
	.datad(tdl_arr_8_11),
	.cin(gnd),
	.combout(\gain_lut_8pts~19_combout ),
	.cout());
defparam \gain_lut_8pts~19 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~20 (
	.dataa(tdl_arr_9_12),
	.datab(tdl_arr_8_12),
	.datac(tdl_arr_9_13),
	.datad(tdl_arr_8_13),
	.cin(gnd),
	.combout(\gain_lut_8pts~20_combout ),
	.cout());
defparam \gain_lut_8pts~20 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~21 (
	.dataa(tdl_arr_9_14),
	.datab(tdl_arr_8_14),
	.datac(tdl_arr_9_15),
	.datad(tdl_arr_8_15),
	.cin(gnd),
	.combout(\gain_lut_8pts~21_combout ),
	.cout());
defparam \gain_lut_8pts~21 .lut_mask = 16'h6996;
defparam \gain_lut_8pts~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~22 (
	.dataa(\gain_lut_8pts~18_combout ),
	.datab(\gain_lut_8pts~19_combout ),
	.datac(\gain_lut_8pts~20_combout ),
	.datad(\gain_lut_8pts~21_combout ),
	.cin(gnd),
	.combout(\gain_lut_8pts~22_combout ),
	.cout());
defparam \gain_lut_8pts~22 .lut_mask = 16'hFFFE;
defparam \gain_lut_8pts~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \gain_lut_8pts~23 (
	.dataa(\gain_lut_8pts~22_combout ),
	.datab(\sdetd.GBLK~q ),
	.datac(\sdetd.ENABLE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\gain_lut_8pts~23_combout ),
	.cout());
defparam \gain_lut_8pts~23 .lut_mask = 16'hFEFE;
defparam \gain_lut_8pts~23 .sum_lutc_input = "datac";

dffeas \gain_lut_8pts[3] (
	.clk(clk),
	.d(\gain_lut_8pts~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_8pts[3]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[3] .is_wysiwyg = "true";
defparam \gain_lut_8pts[3] .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\sdetd.GBLK~q ),
	.datab(\sdetd.ENABLE~q ),
	.datac(\gain_lut_8pts[3]~q ),
	.datad(\gain_lut_blk[3]~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFFFE;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \gain_lut_blk[3] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\gain_lut_blk[3]~q ),
	.prn(vcc));
defparam \gain_lut_blk[3] .is_wysiwyg = "true";
defparam \gain_lut_blk[3] .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\gain_lut_8pts[3]~q ),
	.datab(\gain_lut_blk[3]~q ),
	.datac(gnd),
	.datad(\sdetd.SLBI~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEEFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_rst_1 (
	global_clock_enable,
	tdl_arr_0,
	tdl_arr_01,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	tdl_arr_0;
output 	tdl_arr_01;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~0_combout ;


dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_01),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(tdl_arr_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_cmult_std (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_3_1,
	tdl_arr_3_11,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	clk)/* synthesis synthesis_greybox=1 */;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_5_11;
output 	tdl_arr_9_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_7_1;
output 	tdl_arr_7_11;
output 	tdl_arr_8_1;
output 	tdl_arr_8_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_3_1;
output 	tdl_arr_3_11;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \result_i_tmp[15]~q ;
wire \result_i_tmp[14]~q ;
wire \result_i_tmp[13]~q ;
wire \result_i_tmp[12]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[10]~q ;
wire \result_i_tmp[9]~q ;
wire \result_i_tmp[8]~q ;
wire \result_i_tmp[7]~q ;
wire \result_i_tmp[6]~q ;
wire \result_i_tmp[5]~q ;
wire \result_i_tmp[4]~q ;
wire \result_i_tmp[3]~q ;
wire \result_i_tmp[2]~q ;
wire \result_i_tmp[1]~q ;
wire \result_i_tmp[0]~q ;
wire \result_i_tmp[19]~q ;
wire \result_i_tmp[18]~q ;
wire \result_i_tmp[17]~q ;
wire \result_i_tmp[16]~q ;
wire \result_r_tmp[15]~q ;
wire \result_r_tmp[14]~q ;
wire \result_r_tmp[13]~q ;
wire \result_r_tmp[12]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[10]~q ;
wire \result_r_tmp[9]~q ;
wire \result_r_tmp[8]~q ;
wire \result_r_tmp[7]~q ;
wire \result_r_tmp[6]~q ;
wire \result_r_tmp[5]~q ;
wire \result_r_tmp[4]~q ;
wire \result_r_tmp[3]~q ;
wire \result_r_tmp[2]~q ;
wire \result_r_tmp[1]~q ;
wire \result_r_tmp[0]~q ;
wire \result_r_tmp[19]~q ;
wire \result_r_tmp[18]~q ;
wire \result_r_tmp[17]~q ;
wire \result_r_tmp[16]~q ;


fftsign_asj_fft_tdl \gen_ma:gen_ma_full:imag_delay (
	.data_in({\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_9_1(tdl_arr_9_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_8_1(tdl_arr_8_1),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_3_1(tdl_arr_3_1),
	.clk(clk));

fftsign_asj_fft_tdl_1 \gen_ma:gen_ma_full:real_delay (
	.data_in({\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_9_1(tdl_arr_9_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_8_1(tdl_arr_8_11),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_3_1(tdl_arr_3_11),
	.clk(clk));

fftsign_asj_fft_pround_1 \gen_ma:gen_ma_full:u1 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.result_i_tmp_19(\result_i_tmp[19]~q ),
	.result_i_tmp_18(\result_i_tmp[18]~q ),
	.result_i_tmp_17(\result_i_tmp[17]~q ),
	.result_i_tmp_16(\result_i_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_pround \gen_ma:gen_ma_full:u0 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.result_r_tmp_19(\result_r_tmp[19]~q ),
	.result_r_tmp_18(\result_r_tmp[18]~q ),
	.result_r_tmp_17(\result_r_tmp[17]~q ),
	.result_r_tmp_16(\result_r_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_mult_add \gen_ma:gen_ma_full:ma (
	.dffe5a_15(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.dffe5a_14(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.dffe5a_13(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.dffe5a_12(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.dffe5a_11(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.dffe5a_10(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.dffe5a_9(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.dffe5a_8(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.dffe5a_7(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.dffe5a_6(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.dffe5a_5(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.dffe5a_4(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.dffe5a_3(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.dffe5a_2(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.dffe5a_1(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.dffe5a_0(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.dffe5a_19(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.dffe5a_18(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.dffe5a_17(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.dffe5a_16(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data018(twiddle_data018),
	.twiddle_data019(twiddle_data019),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data008(twiddle_data008),
	.twiddle_data009(twiddle_data009),
	.clk(clk));

fftsign_asj_fft_mult_add_1 \gen_ma:gen_ma_full:ms (
	.dffe7a_15(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.dffe7a_14(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.dffe7a_13(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.dffe7a_12(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.dffe7a_11(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.dffe7a_10(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.dffe7a_9(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.dffe7a_8(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.dffe7a_7(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.dffe7a_6(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.dffe7a_5(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.dffe7a_4(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.dffe7a_3(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.dffe7a_2(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.dffe7a_1(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.dffe7a_0(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.dffe7a_19(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.dffe7a_18(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.dffe7a_17(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.dffe7a_16(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data018(twiddle_data018),
	.twiddle_data019(twiddle_data019),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data008(twiddle_data008),
	.twiddle_data009(twiddle_data009),
	.clk(clk));

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

dffeas \result_i_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[19]~q ),
	.prn(vcc));
defparam \result_i_tmp[19] .is_wysiwyg = "true";
defparam \result_i_tmp[19] .power_up = "low";

dffeas \result_i_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[18]~q ),
	.prn(vcc));
defparam \result_i_tmp[18] .is_wysiwyg = "true";
defparam \result_i_tmp[18] .power_up = "low";

dffeas \result_i_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[17]~q ),
	.prn(vcc));
defparam \result_i_tmp[17] .is_wysiwyg = "true";
defparam \result_i_tmp[17] .power_up = "low";

dffeas \result_i_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[16]~q ),
	.prn(vcc));
defparam \result_i_tmp[16] .is_wysiwyg = "true";
defparam \result_i_tmp[16] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

dffeas \result_r_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[19]~q ),
	.prn(vcc));
defparam \result_r_tmp[19] .is_wysiwyg = "true";
defparam \result_r_tmp[19] .power_up = "low";

dffeas \result_r_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[18]~q ),
	.prn(vcc));
defparam \result_r_tmp[18] .is_wysiwyg = "true";
defparam \result_r_tmp[18] .power_up = "low";

dffeas \result_r_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[17]~q ),
	.prn(vcc));
defparam \result_r_tmp[17] .is_wysiwyg = "true";
defparam \result_r_tmp[17] .power_up = "low";

dffeas \result_r_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[16]~q ),
	.prn(vcc));
defparam \result_r_tmp[16] .is_wysiwyg = "true";
defparam \result_r_tmp[16] .power_up = "low";

endmodule

module fftsign_asj_fft_mult_add (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add MULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data018(twiddle_data018),
	.twiddle_data019(twiddle_data019),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data008(twiddle_data008),
	.twiddle_data009(twiddle_data009),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2,pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,
pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.ena0(global_clock_enable),
	.datab({twiddle_data019,twiddle_data018,twiddle_data017,twiddle_data016,twiddle_data015,twiddle_data014,twiddle_data013,twiddle_data012,twiddle_data011,twiddle_data010,twiddle_data009,twiddle_data008,twiddle_data007,twiddle_data006,twiddle_data005,twiddle_data004,twiddle_data003,
twiddle_data002,twiddle_data001,twiddle_data000}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_1 ALTMULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_1 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_kk6g auto_generated(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_kk6g (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe5a[0]~21 ;
wire \dffe5a[1]~23 ;
wire \dffe5a[2]~25 ;
wire \dffe5a[3]~27 ;
wire \dffe5a[4]~29 ;
wire \dffe5a[5]~31 ;
wire \dffe5a[6]~33 ;
wire \dffe5a[7]~35 ;
wire \dffe5a[8]~37 ;
wire \dffe5a[9]~39 ;
wire \dffe5a[10]~41 ;
wire \dffe5a[11]~43 ;
wire \dffe5a[12]~45 ;
wire \dffe5a[13]~47 ;
wire \dffe5a[14]~49 ;
wire \dffe5a[15]~50_combout ;
wire \dffe5a[14]~48_combout ;
wire \dffe5a[13]~46_combout ;
wire \dffe5a[12]~44_combout ;
wire \dffe5a[11]~42_combout ;
wire \dffe5a[10]~40_combout ;
wire \dffe5a[9]~38_combout ;
wire \dffe5a[8]~36_combout ;
wire \dffe5a[7]~34_combout ;
wire \dffe5a[6]~32_combout ;
wire \dffe5a[5]~30_combout ;
wire \dffe5a[4]~28_combout ;
wire \dffe5a[3]~26_combout ;
wire \dffe5a[2]~24_combout ;
wire \dffe5a[1]~22_combout ;
wire \dffe5a[0]~20_combout ;
wire \dffe5a[15]~51 ;
wire \dffe5a[16]~53 ;
wire \dffe5a[17]~55 ;
wire \dffe5a[18]~57 ;
wire \dffe5a[19]~58_combout ;
wire \dffe5a[18]~56_combout ;
wire \dffe5a[17]~54_combout ;
wire \dffe5a[16]~52_combout ;


fftsign_ded_mult_9a91_1 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe5a[15] (
	.clk(clock0),
	.d(\dffe5a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_15),
	.prn(vcc));
defparam \dffe5a[15] .is_wysiwyg = "true";
defparam \dffe5a[15] .power_up = "low";

dffeas \dffe5a[14] (
	.clk(clock0),
	.d(\dffe5a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_14),
	.prn(vcc));
defparam \dffe5a[14] .is_wysiwyg = "true";
defparam \dffe5a[14] .power_up = "low";

dffeas \dffe5a[13] (
	.clk(clock0),
	.d(\dffe5a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_13),
	.prn(vcc));
defparam \dffe5a[13] .is_wysiwyg = "true";
defparam \dffe5a[13] .power_up = "low";

dffeas \dffe5a[12] (
	.clk(clock0),
	.d(\dffe5a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_12),
	.prn(vcc));
defparam \dffe5a[12] .is_wysiwyg = "true";
defparam \dffe5a[12] .power_up = "low";

dffeas \dffe5a[11] (
	.clk(clock0),
	.d(\dffe5a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_11),
	.prn(vcc));
defparam \dffe5a[11] .is_wysiwyg = "true";
defparam \dffe5a[11] .power_up = "low";

dffeas \dffe5a[10] (
	.clk(clock0),
	.d(\dffe5a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_10),
	.prn(vcc));
defparam \dffe5a[10] .is_wysiwyg = "true";
defparam \dffe5a[10] .power_up = "low";

dffeas \dffe5a[9] (
	.clk(clock0),
	.d(\dffe5a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_9),
	.prn(vcc));
defparam \dffe5a[9] .is_wysiwyg = "true";
defparam \dffe5a[9] .power_up = "low";

dffeas \dffe5a[8] (
	.clk(clock0),
	.d(\dffe5a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_8),
	.prn(vcc));
defparam \dffe5a[8] .is_wysiwyg = "true";
defparam \dffe5a[8] .power_up = "low";

dffeas \dffe5a[7] (
	.clk(clock0),
	.d(\dffe5a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_7),
	.prn(vcc));
defparam \dffe5a[7] .is_wysiwyg = "true";
defparam \dffe5a[7] .power_up = "low";

dffeas \dffe5a[6] (
	.clk(clock0),
	.d(\dffe5a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_6),
	.prn(vcc));
defparam \dffe5a[6] .is_wysiwyg = "true";
defparam \dffe5a[6] .power_up = "low";

dffeas \dffe5a[5] (
	.clk(clock0),
	.d(\dffe5a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_5),
	.prn(vcc));
defparam \dffe5a[5] .is_wysiwyg = "true";
defparam \dffe5a[5] .power_up = "low";

dffeas \dffe5a[4] (
	.clk(clock0),
	.d(\dffe5a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_4),
	.prn(vcc));
defparam \dffe5a[4] .is_wysiwyg = "true";
defparam \dffe5a[4] .power_up = "low";

dffeas \dffe5a[3] (
	.clk(clock0),
	.d(\dffe5a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_3),
	.prn(vcc));
defparam \dffe5a[3] .is_wysiwyg = "true";
defparam \dffe5a[3] .power_up = "low";

dffeas \dffe5a[2] (
	.clk(clock0),
	.d(\dffe5a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_2),
	.prn(vcc));
defparam \dffe5a[2] .is_wysiwyg = "true";
defparam \dffe5a[2] .power_up = "low";

dffeas \dffe5a[1] (
	.clk(clock0),
	.d(\dffe5a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_1),
	.prn(vcc));
defparam \dffe5a[1] .is_wysiwyg = "true";
defparam \dffe5a[1] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock0),
	.d(\dffe5a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_0),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

dffeas \dffe5a[19] (
	.clk(clock0),
	.d(\dffe5a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_19),
	.prn(vcc));
defparam \dffe5a[19] .is_wysiwyg = "true";
defparam \dffe5a[19] .power_up = "low";

dffeas \dffe5a[18] (
	.clk(clock0),
	.d(\dffe5a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_18),
	.prn(vcc));
defparam \dffe5a[18] .is_wysiwyg = "true";
defparam \dffe5a[18] .power_up = "low";

dffeas \dffe5a[17] (
	.clk(clock0),
	.d(\dffe5a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_17),
	.prn(vcc));
defparam \dffe5a[17] .is_wysiwyg = "true";
defparam \dffe5a[17] .power_up = "low";

dffeas \dffe5a[16] (
	.clk(clock0),
	.d(\dffe5a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_16),
	.prn(vcc));
defparam \dffe5a[16] .is_wysiwyg = "true";
defparam \dffe5a[16] .power_up = "low";

cycloneive_lcell_comb \dffe5a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe5a[0]~20_combout ),
	.cout(\dffe5a[0]~21 ));
defparam \dffe5a[0]~20 .lut_mask = 16'h66EE;
defparam \dffe5a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe5a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[0]~21 ),
	.combout(\dffe5a[1]~22_combout ),
	.cout(\dffe5a[1]~23 ));
defparam \dffe5a[1]~22 .lut_mask = 16'h967F;
defparam \dffe5a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[1]~23 ),
	.combout(\dffe5a[2]~24_combout ),
	.cout(\dffe5a[2]~25 ));
defparam \dffe5a[2]~24 .lut_mask = 16'h96EF;
defparam \dffe5a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[2]~25 ),
	.combout(\dffe5a[3]~26_combout ),
	.cout(\dffe5a[3]~27 ));
defparam \dffe5a[3]~26 .lut_mask = 16'h967F;
defparam \dffe5a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[3]~27 ),
	.combout(\dffe5a[4]~28_combout ),
	.cout(\dffe5a[4]~29 ));
defparam \dffe5a[4]~28 .lut_mask = 16'h96EF;
defparam \dffe5a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[4]~29 ),
	.combout(\dffe5a[5]~30_combout ),
	.cout(\dffe5a[5]~31 ));
defparam \dffe5a[5]~30 .lut_mask = 16'h967F;
defparam \dffe5a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[5]~31 ),
	.combout(\dffe5a[6]~32_combout ),
	.cout(\dffe5a[6]~33 ));
defparam \dffe5a[6]~32 .lut_mask = 16'h96EF;
defparam \dffe5a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[6]~33 ),
	.combout(\dffe5a[7]~34_combout ),
	.cout(\dffe5a[7]~35 ));
defparam \dffe5a[7]~34 .lut_mask = 16'h967F;
defparam \dffe5a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[7]~35 ),
	.combout(\dffe5a[8]~36_combout ),
	.cout(\dffe5a[8]~37 ));
defparam \dffe5a[8]~36 .lut_mask = 16'h96EF;
defparam \dffe5a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[8]~37 ),
	.combout(\dffe5a[9]~38_combout ),
	.cout(\dffe5a[9]~39 ));
defparam \dffe5a[9]~38 .lut_mask = 16'h967F;
defparam \dffe5a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[9]~39 ),
	.combout(\dffe5a[10]~40_combout ),
	.cout(\dffe5a[10]~41 ));
defparam \dffe5a[10]~40 .lut_mask = 16'h96EF;
defparam \dffe5a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[10]~41 ),
	.combout(\dffe5a[11]~42_combout ),
	.cout(\dffe5a[11]~43 ));
defparam \dffe5a[11]~42 .lut_mask = 16'h967F;
defparam \dffe5a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[11]~43 ),
	.combout(\dffe5a[12]~44_combout ),
	.cout(\dffe5a[12]~45 ));
defparam \dffe5a[12]~44 .lut_mask = 16'h96EF;
defparam \dffe5a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[12]~45 ),
	.combout(\dffe5a[13]~46_combout ),
	.cout(\dffe5a[13]~47 ));
defparam \dffe5a[13]~46 .lut_mask = 16'h967F;
defparam \dffe5a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[13]~47 ),
	.combout(\dffe5a[14]~48_combout ),
	.cout(\dffe5a[14]~49 ));
defparam \dffe5a[14]~48 .lut_mask = 16'h96EF;
defparam \dffe5a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[14]~49 ),
	.combout(\dffe5a[15]~50_combout ),
	.cout(\dffe5a[15]~51 ));
defparam \dffe5a[15]~50 .lut_mask = 16'h967F;
defparam \dffe5a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[15]~51 ),
	.combout(\dffe5a[16]~52_combout ),
	.cout(\dffe5a[16]~53 ));
defparam \dffe5a[16]~52 .lut_mask = 16'h96EF;
defparam \dffe5a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[16]~53 ),
	.combout(\dffe5a[17]~54_combout ),
	.cout(\dffe5a[17]~55 ));
defparam \dffe5a[17]~54 .lut_mask = 16'h967F;
defparam \dffe5a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[17]~55 ),
	.combout(\dffe5a[18]~56_combout ),
	.cout(\dffe5a[18]~57 ));
defparam \dffe5a[18]~56 .lut_mask = 16'h96EF;
defparam \dffe5a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe5a[18]~57 ),
	.combout(\dffe5a[19]~58_combout ),
	.cout());
defparam \dffe5a[19]~58 .lut_mask = 16'h9696;
defparam \dffe5a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_1 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_mult_add_1 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_1 MULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data018(twiddle_data018),
	.twiddle_data019(twiddle_data019),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.twiddle_data007(twiddle_data007),
	.twiddle_data008(twiddle_data008),
	.twiddle_data009(twiddle_data009),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add_1 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data018,
	twiddle_data019,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data007,
	twiddle_data008,
	twiddle_data009,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data018;
input 	twiddle_data019;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data007;
input 	twiddle_data008;
input 	twiddle_data009;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old_1 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21,pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,
pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.ena0(global_clock_enable),
	.datab({twiddle_data019,twiddle_data018,twiddle_data017,twiddle_data016,twiddle_data015,twiddle_data014,twiddle_data013,twiddle_data012,twiddle_data011,twiddle_data010,twiddle_data009,twiddle_data008,twiddle_data007,twiddle_data006,twiddle_data005,twiddle_data004,twiddle_data003,
twiddle_data002,twiddle_data001,twiddle_data000}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old_1 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_2 ALTMULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_2 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_ll6g auto_generated(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_ll6g (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe7a[0]~21 ;
wire \dffe7a[1]~23 ;
wire \dffe7a[2]~25 ;
wire \dffe7a[3]~27 ;
wire \dffe7a[4]~29 ;
wire \dffe7a[5]~31 ;
wire \dffe7a[6]~33 ;
wire \dffe7a[7]~35 ;
wire \dffe7a[8]~37 ;
wire \dffe7a[9]~39 ;
wire \dffe7a[10]~41 ;
wire \dffe7a[11]~43 ;
wire \dffe7a[12]~45 ;
wire \dffe7a[13]~47 ;
wire \dffe7a[14]~49 ;
wire \dffe7a[15]~50_combout ;
wire \dffe7a[14]~48_combout ;
wire \dffe7a[13]~46_combout ;
wire \dffe7a[12]~44_combout ;
wire \dffe7a[11]~42_combout ;
wire \dffe7a[10]~40_combout ;
wire \dffe7a[9]~38_combout ;
wire \dffe7a[8]~36_combout ;
wire \dffe7a[7]~34_combout ;
wire \dffe7a[6]~32_combout ;
wire \dffe7a[5]~30_combout ;
wire \dffe7a[4]~28_combout ;
wire \dffe7a[3]~26_combout ;
wire \dffe7a[2]~24_combout ;
wire \dffe7a[1]~22_combout ;
wire \dffe7a[0]~20_combout ;
wire \dffe7a[15]~51 ;
wire \dffe7a[16]~53 ;
wire \dffe7a[17]~55 ;
wire \dffe7a[18]~57 ;
wire \dffe7a[19]~58_combout ;
wire \dffe7a[18]~56_combout ;
wire \dffe7a[17]~54_combout ;
wire \dffe7a[16]~52_combout ;


fftsign_ded_mult_9a91_3 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91_2 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe7a[15] (
	.clk(clock0),
	.d(\dffe7a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_15),
	.prn(vcc));
defparam \dffe7a[15] .is_wysiwyg = "true";
defparam \dffe7a[15] .power_up = "low";

dffeas \dffe7a[14] (
	.clk(clock0),
	.d(\dffe7a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_14),
	.prn(vcc));
defparam \dffe7a[14] .is_wysiwyg = "true";
defparam \dffe7a[14] .power_up = "low";

dffeas \dffe7a[13] (
	.clk(clock0),
	.d(\dffe7a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_13),
	.prn(vcc));
defparam \dffe7a[13] .is_wysiwyg = "true";
defparam \dffe7a[13] .power_up = "low";

dffeas \dffe7a[12] (
	.clk(clock0),
	.d(\dffe7a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_12),
	.prn(vcc));
defparam \dffe7a[12] .is_wysiwyg = "true";
defparam \dffe7a[12] .power_up = "low";

dffeas \dffe7a[11] (
	.clk(clock0),
	.d(\dffe7a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_11),
	.prn(vcc));
defparam \dffe7a[11] .is_wysiwyg = "true";
defparam \dffe7a[11] .power_up = "low";

dffeas \dffe7a[10] (
	.clk(clock0),
	.d(\dffe7a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_10),
	.prn(vcc));
defparam \dffe7a[10] .is_wysiwyg = "true";
defparam \dffe7a[10] .power_up = "low";

dffeas \dffe7a[9] (
	.clk(clock0),
	.d(\dffe7a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_9),
	.prn(vcc));
defparam \dffe7a[9] .is_wysiwyg = "true";
defparam \dffe7a[9] .power_up = "low";

dffeas \dffe7a[8] (
	.clk(clock0),
	.d(\dffe7a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_8),
	.prn(vcc));
defparam \dffe7a[8] .is_wysiwyg = "true";
defparam \dffe7a[8] .power_up = "low";

dffeas \dffe7a[7] (
	.clk(clock0),
	.d(\dffe7a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_7),
	.prn(vcc));
defparam \dffe7a[7] .is_wysiwyg = "true";
defparam \dffe7a[7] .power_up = "low";

dffeas \dffe7a[6] (
	.clk(clock0),
	.d(\dffe7a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_6),
	.prn(vcc));
defparam \dffe7a[6] .is_wysiwyg = "true";
defparam \dffe7a[6] .power_up = "low";

dffeas \dffe7a[5] (
	.clk(clock0),
	.d(\dffe7a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_5),
	.prn(vcc));
defparam \dffe7a[5] .is_wysiwyg = "true";
defparam \dffe7a[5] .power_up = "low";

dffeas \dffe7a[4] (
	.clk(clock0),
	.d(\dffe7a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_4),
	.prn(vcc));
defparam \dffe7a[4] .is_wysiwyg = "true";
defparam \dffe7a[4] .power_up = "low";

dffeas \dffe7a[3] (
	.clk(clock0),
	.d(\dffe7a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_3),
	.prn(vcc));
defparam \dffe7a[3] .is_wysiwyg = "true";
defparam \dffe7a[3] .power_up = "low";

dffeas \dffe7a[2] (
	.clk(clock0),
	.d(\dffe7a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_2),
	.prn(vcc));
defparam \dffe7a[2] .is_wysiwyg = "true";
defparam \dffe7a[2] .power_up = "low";

dffeas \dffe7a[1] (
	.clk(clock0),
	.d(\dffe7a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_1),
	.prn(vcc));
defparam \dffe7a[1] .is_wysiwyg = "true";
defparam \dffe7a[1] .power_up = "low";

dffeas \dffe7a[0] (
	.clk(clock0),
	.d(\dffe7a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_0),
	.prn(vcc));
defparam \dffe7a[0] .is_wysiwyg = "true";
defparam \dffe7a[0] .power_up = "low";

dffeas \dffe7a[19] (
	.clk(clock0),
	.d(\dffe7a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_19),
	.prn(vcc));
defparam \dffe7a[19] .is_wysiwyg = "true";
defparam \dffe7a[19] .power_up = "low";

dffeas \dffe7a[18] (
	.clk(clock0),
	.d(\dffe7a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_18),
	.prn(vcc));
defparam \dffe7a[18] .is_wysiwyg = "true";
defparam \dffe7a[18] .power_up = "low";

dffeas \dffe7a[17] (
	.clk(clock0),
	.d(\dffe7a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_17),
	.prn(vcc));
defparam \dffe7a[17] .is_wysiwyg = "true";
defparam \dffe7a[17] .power_up = "low";

dffeas \dffe7a[16] (
	.clk(clock0),
	.d(\dffe7a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_16),
	.prn(vcc));
defparam \dffe7a[16] .is_wysiwyg = "true";
defparam \dffe7a[16] .power_up = "low";

cycloneive_lcell_comb \dffe7a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe7a[0]~20_combout ),
	.cout(\dffe7a[0]~21 ));
defparam \dffe7a[0]~20 .lut_mask = 16'h66DD;
defparam \dffe7a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe7a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[0]~21 ),
	.combout(\dffe7a[1]~22_combout ),
	.cout(\dffe7a[1]~23 ));
defparam \dffe7a[1]~22 .lut_mask = 16'h96BF;
defparam \dffe7a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[1]~23 ),
	.combout(\dffe7a[2]~24_combout ),
	.cout(\dffe7a[2]~25 ));
defparam \dffe7a[2]~24 .lut_mask = 16'h96DF;
defparam \dffe7a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[2]~25 ),
	.combout(\dffe7a[3]~26_combout ),
	.cout(\dffe7a[3]~27 ));
defparam \dffe7a[3]~26 .lut_mask = 16'h96BF;
defparam \dffe7a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[3]~27 ),
	.combout(\dffe7a[4]~28_combout ),
	.cout(\dffe7a[4]~29 ));
defparam \dffe7a[4]~28 .lut_mask = 16'h96DF;
defparam \dffe7a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[4]~29 ),
	.combout(\dffe7a[5]~30_combout ),
	.cout(\dffe7a[5]~31 ));
defparam \dffe7a[5]~30 .lut_mask = 16'h96BF;
defparam \dffe7a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[5]~31 ),
	.combout(\dffe7a[6]~32_combout ),
	.cout(\dffe7a[6]~33 ));
defparam \dffe7a[6]~32 .lut_mask = 16'h96DF;
defparam \dffe7a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[6]~33 ),
	.combout(\dffe7a[7]~34_combout ),
	.cout(\dffe7a[7]~35 ));
defparam \dffe7a[7]~34 .lut_mask = 16'h96BF;
defparam \dffe7a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[7]~35 ),
	.combout(\dffe7a[8]~36_combout ),
	.cout(\dffe7a[8]~37 ));
defparam \dffe7a[8]~36 .lut_mask = 16'h96DF;
defparam \dffe7a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[8]~37 ),
	.combout(\dffe7a[9]~38_combout ),
	.cout(\dffe7a[9]~39 ));
defparam \dffe7a[9]~38 .lut_mask = 16'h96BF;
defparam \dffe7a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[9]~39 ),
	.combout(\dffe7a[10]~40_combout ),
	.cout(\dffe7a[10]~41 ));
defparam \dffe7a[10]~40 .lut_mask = 16'h96DF;
defparam \dffe7a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[10]~41 ),
	.combout(\dffe7a[11]~42_combout ),
	.cout(\dffe7a[11]~43 ));
defparam \dffe7a[11]~42 .lut_mask = 16'h96BF;
defparam \dffe7a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[11]~43 ),
	.combout(\dffe7a[12]~44_combout ),
	.cout(\dffe7a[12]~45 ));
defparam \dffe7a[12]~44 .lut_mask = 16'h96DF;
defparam \dffe7a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[12]~45 ),
	.combout(\dffe7a[13]~46_combout ),
	.cout(\dffe7a[13]~47 ));
defparam \dffe7a[13]~46 .lut_mask = 16'h96BF;
defparam \dffe7a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[13]~47 ),
	.combout(\dffe7a[14]~48_combout ),
	.cout(\dffe7a[14]~49 ));
defparam \dffe7a[14]~48 .lut_mask = 16'h96DF;
defparam \dffe7a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[14]~49 ),
	.combout(\dffe7a[15]~50_combout ),
	.cout(\dffe7a[15]~51 ));
defparam \dffe7a[15]~50 .lut_mask = 16'h96BF;
defparam \dffe7a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[15]~51 ),
	.combout(\dffe7a[16]~52_combout ),
	.cout(\dffe7a[16]~53 ));
defparam \dffe7a[16]~52 .lut_mask = 16'h96DF;
defparam \dffe7a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[16]~53 ),
	.combout(\dffe7a[17]~54_combout ),
	.cout(\dffe7a[17]~55 ));
defparam \dffe7a[17]~54 .lut_mask = 16'h96BF;
defparam \dffe7a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[17]~55 ),
	.combout(\dffe7a[18]~56_combout ),
	.cout(\dffe7a[18]~57 ));
defparam \dffe7a[18]~56 .lut_mask = 16'h96DF;
defparam \dffe7a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe7a[18]~57 ),
	.combout(\dffe7a[19]~58_combout ),
	.cout());
defparam \dffe7a[19]~58 .lut_mask = 16'h9696;
defparam \dffe7a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91_2 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_3 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_pround (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_1 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_1 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_r_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_r_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_r_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_r_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_r_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_r_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_r_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_r_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_r_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_r_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_r_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_r_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_r_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_r_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_r_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_r_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_r_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_r_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_r_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_1 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_2 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_2 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj_1 auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj_1 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_i_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_i_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_i_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_i_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_i_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_i_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_i_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_i_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_i_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_i_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_i_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_i_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_i_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_i_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_i_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_i_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_i_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_i_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_i_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm1|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_tdl (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_tdl_1 (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_cmult_std_1 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_3_1,
	tdl_arr_3_11,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	clk)/* synthesis synthesis_greybox=1 */;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_5_11;
output 	tdl_arr_9_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_7_1;
output 	tdl_arr_7_11;
output 	tdl_arr_8_1;
output 	tdl_arr_8_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_3_1;
output 	tdl_arr_3_11;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \result_i_tmp[15]~q ;
wire \result_i_tmp[14]~q ;
wire \result_i_tmp[13]~q ;
wire \result_i_tmp[12]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[10]~q ;
wire \result_i_tmp[9]~q ;
wire \result_i_tmp[8]~q ;
wire \result_i_tmp[7]~q ;
wire \result_i_tmp[6]~q ;
wire \result_i_tmp[5]~q ;
wire \result_i_tmp[4]~q ;
wire \result_i_tmp[3]~q ;
wire \result_i_tmp[2]~q ;
wire \result_i_tmp[1]~q ;
wire \result_i_tmp[0]~q ;
wire \result_i_tmp[19]~q ;
wire \result_i_tmp[18]~q ;
wire \result_i_tmp[17]~q ;
wire \result_i_tmp[16]~q ;
wire \result_r_tmp[15]~q ;
wire \result_r_tmp[14]~q ;
wire \result_r_tmp[13]~q ;
wire \result_r_tmp[12]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[10]~q ;
wire \result_r_tmp[9]~q ;
wire \result_r_tmp[8]~q ;
wire \result_r_tmp[7]~q ;
wire \result_r_tmp[6]~q ;
wire \result_r_tmp[5]~q ;
wire \result_r_tmp[4]~q ;
wire \result_r_tmp[3]~q ;
wire \result_r_tmp[2]~q ;
wire \result_r_tmp[1]~q ;
wire \result_r_tmp[0]~q ;
wire \result_r_tmp[19]~q ;
wire \result_r_tmp[18]~q ;
wire \result_r_tmp[17]~q ;
wire \result_r_tmp[16]~q ;


fftsign_asj_fft_tdl_2 \gen_ma:gen_ma_full:imag_delay (
	.data_in({\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_9_1(tdl_arr_9_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_8_1(tdl_arr_8_1),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_3_1(tdl_arr_3_1),
	.clk(clk));

fftsign_asj_fft_tdl_3 \gen_ma:gen_ma_full:real_delay (
	.data_in({\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_9_1(tdl_arr_9_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_8_1(tdl_arr_8_11),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_3_1(tdl_arr_3_11),
	.clk(clk));

fftsign_asj_fft_pround_3 \gen_ma:gen_ma_full:u1 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.result_i_tmp_19(\result_i_tmp[19]~q ),
	.result_i_tmp_18(\result_i_tmp[18]~q ),
	.result_i_tmp_17(\result_i_tmp[17]~q ),
	.result_i_tmp_16(\result_i_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_pround_2 \gen_ma:gen_ma_full:u0 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.result_r_tmp_19(\result_r_tmp[19]~q ),
	.result_r_tmp_18(\result_r_tmp[18]~q ),
	.result_r_tmp_17(\result_r_tmp[17]~q ),
	.result_r_tmp_16(\result_r_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_mult_add_2 \gen_ma:gen_ma_full:ma (
	.dffe5a_15(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.dffe5a_14(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.dffe5a_13(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.dffe5a_12(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.dffe5a_11(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.dffe5a_10(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.dffe5a_9(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.dffe5a_8(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.dffe5a_7(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.dffe5a_6(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.dffe5a_5(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.dffe5a_4(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.dffe5a_3(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.dffe5a_2(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.dffe5a_1(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.dffe5a_0(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.dffe5a_19(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.dffe5a_18(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.dffe5a_17(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.dffe5a_16(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.twiddle_data118(twiddle_data118),
	.twiddle_data119(twiddle_data119),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data108(twiddle_data108),
	.twiddle_data109(twiddle_data109),
	.clk(clk));

fftsign_asj_fft_mult_add_3 \gen_ma:gen_ma_full:ms (
	.dffe7a_15(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.dffe7a_14(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.dffe7a_13(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.dffe7a_12(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.dffe7a_11(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.dffe7a_10(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.dffe7a_9(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.dffe7a_8(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.dffe7a_7(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.dffe7a_6(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.dffe7a_5(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.dffe7a_4(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.dffe7a_3(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.dffe7a_2(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.dffe7a_1(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.dffe7a_0(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.dffe7a_19(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.dffe7a_18(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.dffe7a_17(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.dffe7a_16(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.twiddle_data118(twiddle_data118),
	.twiddle_data119(twiddle_data119),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data108(twiddle_data108),
	.twiddle_data109(twiddle_data109),
	.clk(clk));

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

dffeas \result_i_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[19]~q ),
	.prn(vcc));
defparam \result_i_tmp[19] .is_wysiwyg = "true";
defparam \result_i_tmp[19] .power_up = "low";

dffeas \result_i_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[18]~q ),
	.prn(vcc));
defparam \result_i_tmp[18] .is_wysiwyg = "true";
defparam \result_i_tmp[18] .power_up = "low";

dffeas \result_i_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[17]~q ),
	.prn(vcc));
defparam \result_i_tmp[17] .is_wysiwyg = "true";
defparam \result_i_tmp[17] .power_up = "low";

dffeas \result_i_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[16]~q ),
	.prn(vcc));
defparam \result_i_tmp[16] .is_wysiwyg = "true";
defparam \result_i_tmp[16] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

dffeas \result_r_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[19]~q ),
	.prn(vcc));
defparam \result_r_tmp[19] .is_wysiwyg = "true";
defparam \result_r_tmp[19] .power_up = "low";

dffeas \result_r_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[18]~q ),
	.prn(vcc));
defparam \result_r_tmp[18] .is_wysiwyg = "true";
defparam \result_r_tmp[18] .power_up = "low";

dffeas \result_r_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[17]~q ),
	.prn(vcc));
defparam \result_r_tmp[17] .is_wysiwyg = "true";
defparam \result_r_tmp[17] .power_up = "low";

dffeas \result_r_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[16]~q ),
	.prn(vcc));
defparam \result_r_tmp[16] .is_wysiwyg = "true";
defparam \result_r_tmp[16] .power_up = "low";

endmodule

module fftsign_asj_fft_mult_add_2 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_2 MULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.twiddle_data118(twiddle_data118),
	.twiddle_data119(twiddle_data119),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data108(twiddle_data108),
	.twiddle_data109(twiddle_data109),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add_2 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old_2 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2,pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,
pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.ena0(global_clock_enable),
	.datab({twiddle_data119,twiddle_data118,twiddle_data117,twiddle_data116,twiddle_data115,twiddle_data114,twiddle_data113,twiddle_data112,twiddle_data111,twiddle_data110,twiddle_data109,twiddle_data108,twiddle_data107,twiddle_data106,twiddle_data105,twiddle_data104,twiddle_data103,
twiddle_data102,twiddle_data101,twiddle_data100}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old_2 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_3 ALTMULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_3 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_kk6g_1 auto_generated(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_kk6g_1 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe5a[0]~21 ;
wire \dffe5a[1]~23 ;
wire \dffe5a[2]~25 ;
wire \dffe5a[3]~27 ;
wire \dffe5a[4]~29 ;
wire \dffe5a[5]~31 ;
wire \dffe5a[6]~33 ;
wire \dffe5a[7]~35 ;
wire \dffe5a[8]~37 ;
wire \dffe5a[9]~39 ;
wire \dffe5a[10]~41 ;
wire \dffe5a[11]~43 ;
wire \dffe5a[12]~45 ;
wire \dffe5a[13]~47 ;
wire \dffe5a[14]~49 ;
wire \dffe5a[15]~50_combout ;
wire \dffe5a[14]~48_combout ;
wire \dffe5a[13]~46_combout ;
wire \dffe5a[12]~44_combout ;
wire \dffe5a[11]~42_combout ;
wire \dffe5a[10]~40_combout ;
wire \dffe5a[9]~38_combout ;
wire \dffe5a[8]~36_combout ;
wire \dffe5a[7]~34_combout ;
wire \dffe5a[6]~32_combout ;
wire \dffe5a[5]~30_combout ;
wire \dffe5a[4]~28_combout ;
wire \dffe5a[3]~26_combout ;
wire \dffe5a[2]~24_combout ;
wire \dffe5a[1]~22_combout ;
wire \dffe5a[0]~20_combout ;
wire \dffe5a[15]~51 ;
wire \dffe5a[16]~53 ;
wire \dffe5a[17]~55 ;
wire \dffe5a[18]~57 ;
wire \dffe5a[19]~58_combout ;
wire \dffe5a[18]~56_combout ;
wire \dffe5a[17]~54_combout ;
wire \dffe5a[16]~52_combout ;


fftsign_ded_mult_9a91_5 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91_4 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe5a[15] (
	.clk(clock0),
	.d(\dffe5a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_15),
	.prn(vcc));
defparam \dffe5a[15] .is_wysiwyg = "true";
defparam \dffe5a[15] .power_up = "low";

dffeas \dffe5a[14] (
	.clk(clock0),
	.d(\dffe5a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_14),
	.prn(vcc));
defparam \dffe5a[14] .is_wysiwyg = "true";
defparam \dffe5a[14] .power_up = "low";

dffeas \dffe5a[13] (
	.clk(clock0),
	.d(\dffe5a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_13),
	.prn(vcc));
defparam \dffe5a[13] .is_wysiwyg = "true";
defparam \dffe5a[13] .power_up = "low";

dffeas \dffe5a[12] (
	.clk(clock0),
	.d(\dffe5a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_12),
	.prn(vcc));
defparam \dffe5a[12] .is_wysiwyg = "true";
defparam \dffe5a[12] .power_up = "low";

dffeas \dffe5a[11] (
	.clk(clock0),
	.d(\dffe5a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_11),
	.prn(vcc));
defparam \dffe5a[11] .is_wysiwyg = "true";
defparam \dffe5a[11] .power_up = "low";

dffeas \dffe5a[10] (
	.clk(clock0),
	.d(\dffe5a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_10),
	.prn(vcc));
defparam \dffe5a[10] .is_wysiwyg = "true";
defparam \dffe5a[10] .power_up = "low";

dffeas \dffe5a[9] (
	.clk(clock0),
	.d(\dffe5a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_9),
	.prn(vcc));
defparam \dffe5a[9] .is_wysiwyg = "true";
defparam \dffe5a[9] .power_up = "low";

dffeas \dffe5a[8] (
	.clk(clock0),
	.d(\dffe5a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_8),
	.prn(vcc));
defparam \dffe5a[8] .is_wysiwyg = "true";
defparam \dffe5a[8] .power_up = "low";

dffeas \dffe5a[7] (
	.clk(clock0),
	.d(\dffe5a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_7),
	.prn(vcc));
defparam \dffe5a[7] .is_wysiwyg = "true";
defparam \dffe5a[7] .power_up = "low";

dffeas \dffe5a[6] (
	.clk(clock0),
	.d(\dffe5a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_6),
	.prn(vcc));
defparam \dffe5a[6] .is_wysiwyg = "true";
defparam \dffe5a[6] .power_up = "low";

dffeas \dffe5a[5] (
	.clk(clock0),
	.d(\dffe5a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_5),
	.prn(vcc));
defparam \dffe5a[5] .is_wysiwyg = "true";
defparam \dffe5a[5] .power_up = "low";

dffeas \dffe5a[4] (
	.clk(clock0),
	.d(\dffe5a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_4),
	.prn(vcc));
defparam \dffe5a[4] .is_wysiwyg = "true";
defparam \dffe5a[4] .power_up = "low";

dffeas \dffe5a[3] (
	.clk(clock0),
	.d(\dffe5a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_3),
	.prn(vcc));
defparam \dffe5a[3] .is_wysiwyg = "true";
defparam \dffe5a[3] .power_up = "low";

dffeas \dffe5a[2] (
	.clk(clock0),
	.d(\dffe5a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_2),
	.prn(vcc));
defparam \dffe5a[2] .is_wysiwyg = "true";
defparam \dffe5a[2] .power_up = "low";

dffeas \dffe5a[1] (
	.clk(clock0),
	.d(\dffe5a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_1),
	.prn(vcc));
defparam \dffe5a[1] .is_wysiwyg = "true";
defparam \dffe5a[1] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock0),
	.d(\dffe5a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_0),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

dffeas \dffe5a[19] (
	.clk(clock0),
	.d(\dffe5a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_19),
	.prn(vcc));
defparam \dffe5a[19] .is_wysiwyg = "true";
defparam \dffe5a[19] .power_up = "low";

dffeas \dffe5a[18] (
	.clk(clock0),
	.d(\dffe5a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_18),
	.prn(vcc));
defparam \dffe5a[18] .is_wysiwyg = "true";
defparam \dffe5a[18] .power_up = "low";

dffeas \dffe5a[17] (
	.clk(clock0),
	.d(\dffe5a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_17),
	.prn(vcc));
defparam \dffe5a[17] .is_wysiwyg = "true";
defparam \dffe5a[17] .power_up = "low";

dffeas \dffe5a[16] (
	.clk(clock0),
	.d(\dffe5a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_16),
	.prn(vcc));
defparam \dffe5a[16] .is_wysiwyg = "true";
defparam \dffe5a[16] .power_up = "low";

cycloneive_lcell_comb \dffe5a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe5a[0]~20_combout ),
	.cout(\dffe5a[0]~21 ));
defparam \dffe5a[0]~20 .lut_mask = 16'h66EE;
defparam \dffe5a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe5a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[0]~21 ),
	.combout(\dffe5a[1]~22_combout ),
	.cout(\dffe5a[1]~23 ));
defparam \dffe5a[1]~22 .lut_mask = 16'h967F;
defparam \dffe5a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[1]~23 ),
	.combout(\dffe5a[2]~24_combout ),
	.cout(\dffe5a[2]~25 ));
defparam \dffe5a[2]~24 .lut_mask = 16'h96EF;
defparam \dffe5a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[2]~25 ),
	.combout(\dffe5a[3]~26_combout ),
	.cout(\dffe5a[3]~27 ));
defparam \dffe5a[3]~26 .lut_mask = 16'h967F;
defparam \dffe5a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[3]~27 ),
	.combout(\dffe5a[4]~28_combout ),
	.cout(\dffe5a[4]~29 ));
defparam \dffe5a[4]~28 .lut_mask = 16'h96EF;
defparam \dffe5a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[4]~29 ),
	.combout(\dffe5a[5]~30_combout ),
	.cout(\dffe5a[5]~31 ));
defparam \dffe5a[5]~30 .lut_mask = 16'h967F;
defparam \dffe5a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[5]~31 ),
	.combout(\dffe5a[6]~32_combout ),
	.cout(\dffe5a[6]~33 ));
defparam \dffe5a[6]~32 .lut_mask = 16'h96EF;
defparam \dffe5a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[6]~33 ),
	.combout(\dffe5a[7]~34_combout ),
	.cout(\dffe5a[7]~35 ));
defparam \dffe5a[7]~34 .lut_mask = 16'h967F;
defparam \dffe5a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[7]~35 ),
	.combout(\dffe5a[8]~36_combout ),
	.cout(\dffe5a[8]~37 ));
defparam \dffe5a[8]~36 .lut_mask = 16'h96EF;
defparam \dffe5a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[8]~37 ),
	.combout(\dffe5a[9]~38_combout ),
	.cout(\dffe5a[9]~39 ));
defparam \dffe5a[9]~38 .lut_mask = 16'h967F;
defparam \dffe5a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[9]~39 ),
	.combout(\dffe5a[10]~40_combout ),
	.cout(\dffe5a[10]~41 ));
defparam \dffe5a[10]~40 .lut_mask = 16'h96EF;
defparam \dffe5a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[10]~41 ),
	.combout(\dffe5a[11]~42_combout ),
	.cout(\dffe5a[11]~43 ));
defparam \dffe5a[11]~42 .lut_mask = 16'h967F;
defparam \dffe5a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[11]~43 ),
	.combout(\dffe5a[12]~44_combout ),
	.cout(\dffe5a[12]~45 ));
defparam \dffe5a[12]~44 .lut_mask = 16'h96EF;
defparam \dffe5a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[12]~45 ),
	.combout(\dffe5a[13]~46_combout ),
	.cout(\dffe5a[13]~47 ));
defparam \dffe5a[13]~46 .lut_mask = 16'h967F;
defparam \dffe5a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[13]~47 ),
	.combout(\dffe5a[14]~48_combout ),
	.cout(\dffe5a[14]~49 ));
defparam \dffe5a[14]~48 .lut_mask = 16'h96EF;
defparam \dffe5a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[14]~49 ),
	.combout(\dffe5a[15]~50_combout ),
	.cout(\dffe5a[15]~51 ));
defparam \dffe5a[15]~50 .lut_mask = 16'h967F;
defparam \dffe5a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[15]~51 ),
	.combout(\dffe5a[16]~52_combout ),
	.cout(\dffe5a[16]~53 ));
defparam \dffe5a[16]~52 .lut_mask = 16'h96EF;
defparam \dffe5a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[16]~53 ),
	.combout(\dffe5a[17]~54_combout ),
	.cout(\dffe5a[17]~55 ));
defparam \dffe5a[17]~54 .lut_mask = 16'h967F;
defparam \dffe5a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[17]~55 ),
	.combout(\dffe5a[18]~56_combout ),
	.cout(\dffe5a[18]~57 ));
defparam \dffe5a[18]~56 .lut_mask = 16'h96EF;
defparam \dffe5a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe5a[18]~57 ),
	.combout(\dffe5a[19]~58_combout ),
	.cout());
defparam \dffe5a[19]~58 .lut_mask = 16'h9696;
defparam \dffe5a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91_4 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_5 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_mult_add_3 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_3 MULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.twiddle_data118(twiddle_data118),
	.twiddle_data119(twiddle_data119),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.twiddle_data107(twiddle_data107),
	.twiddle_data108(twiddle_data108),
	.twiddle_data109(twiddle_data109),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add_3 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data118,
	twiddle_data119,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data107,
	twiddle_data108,
	twiddle_data109,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data118;
input 	twiddle_data119;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data107;
input 	twiddle_data108;
input 	twiddle_data109;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old_3 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21,pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,
pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.ena0(global_clock_enable),
	.datab({twiddle_data119,twiddle_data118,twiddle_data117,twiddle_data116,twiddle_data115,twiddle_data114,twiddle_data113,twiddle_data112,twiddle_data111,twiddle_data110,twiddle_data109,twiddle_data108,twiddle_data107,twiddle_data106,twiddle_data105,twiddle_data104,twiddle_data103,
twiddle_data102,twiddle_data101,twiddle_data100}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old_3 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_4 ALTMULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_4 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_ll6g_1 auto_generated(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_ll6g_1 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe7a[0]~21 ;
wire \dffe7a[1]~23 ;
wire \dffe7a[2]~25 ;
wire \dffe7a[3]~27 ;
wire \dffe7a[4]~29 ;
wire \dffe7a[5]~31 ;
wire \dffe7a[6]~33 ;
wire \dffe7a[7]~35 ;
wire \dffe7a[8]~37 ;
wire \dffe7a[9]~39 ;
wire \dffe7a[10]~41 ;
wire \dffe7a[11]~43 ;
wire \dffe7a[12]~45 ;
wire \dffe7a[13]~47 ;
wire \dffe7a[14]~49 ;
wire \dffe7a[15]~50_combout ;
wire \dffe7a[14]~48_combout ;
wire \dffe7a[13]~46_combout ;
wire \dffe7a[12]~44_combout ;
wire \dffe7a[11]~42_combout ;
wire \dffe7a[10]~40_combout ;
wire \dffe7a[9]~38_combout ;
wire \dffe7a[8]~36_combout ;
wire \dffe7a[7]~34_combout ;
wire \dffe7a[6]~32_combout ;
wire \dffe7a[5]~30_combout ;
wire \dffe7a[4]~28_combout ;
wire \dffe7a[3]~26_combout ;
wire \dffe7a[2]~24_combout ;
wire \dffe7a[1]~22_combout ;
wire \dffe7a[0]~20_combout ;
wire \dffe7a[15]~51 ;
wire \dffe7a[16]~53 ;
wire \dffe7a[17]~55 ;
wire \dffe7a[18]~57 ;
wire \dffe7a[19]~58_combout ;
wire \dffe7a[18]~56_combout ;
wire \dffe7a[17]~54_combout ;
wire \dffe7a[16]~52_combout ;


fftsign_ded_mult_9a91_7 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91_6 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe7a[15] (
	.clk(clock0),
	.d(\dffe7a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_15),
	.prn(vcc));
defparam \dffe7a[15] .is_wysiwyg = "true";
defparam \dffe7a[15] .power_up = "low";

dffeas \dffe7a[14] (
	.clk(clock0),
	.d(\dffe7a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_14),
	.prn(vcc));
defparam \dffe7a[14] .is_wysiwyg = "true";
defparam \dffe7a[14] .power_up = "low";

dffeas \dffe7a[13] (
	.clk(clock0),
	.d(\dffe7a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_13),
	.prn(vcc));
defparam \dffe7a[13] .is_wysiwyg = "true";
defparam \dffe7a[13] .power_up = "low";

dffeas \dffe7a[12] (
	.clk(clock0),
	.d(\dffe7a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_12),
	.prn(vcc));
defparam \dffe7a[12] .is_wysiwyg = "true";
defparam \dffe7a[12] .power_up = "low";

dffeas \dffe7a[11] (
	.clk(clock0),
	.d(\dffe7a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_11),
	.prn(vcc));
defparam \dffe7a[11] .is_wysiwyg = "true";
defparam \dffe7a[11] .power_up = "low";

dffeas \dffe7a[10] (
	.clk(clock0),
	.d(\dffe7a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_10),
	.prn(vcc));
defparam \dffe7a[10] .is_wysiwyg = "true";
defparam \dffe7a[10] .power_up = "low";

dffeas \dffe7a[9] (
	.clk(clock0),
	.d(\dffe7a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_9),
	.prn(vcc));
defparam \dffe7a[9] .is_wysiwyg = "true";
defparam \dffe7a[9] .power_up = "low";

dffeas \dffe7a[8] (
	.clk(clock0),
	.d(\dffe7a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_8),
	.prn(vcc));
defparam \dffe7a[8] .is_wysiwyg = "true";
defparam \dffe7a[8] .power_up = "low";

dffeas \dffe7a[7] (
	.clk(clock0),
	.d(\dffe7a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_7),
	.prn(vcc));
defparam \dffe7a[7] .is_wysiwyg = "true";
defparam \dffe7a[7] .power_up = "low";

dffeas \dffe7a[6] (
	.clk(clock0),
	.d(\dffe7a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_6),
	.prn(vcc));
defparam \dffe7a[6] .is_wysiwyg = "true";
defparam \dffe7a[6] .power_up = "low";

dffeas \dffe7a[5] (
	.clk(clock0),
	.d(\dffe7a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_5),
	.prn(vcc));
defparam \dffe7a[5] .is_wysiwyg = "true";
defparam \dffe7a[5] .power_up = "low";

dffeas \dffe7a[4] (
	.clk(clock0),
	.d(\dffe7a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_4),
	.prn(vcc));
defparam \dffe7a[4] .is_wysiwyg = "true";
defparam \dffe7a[4] .power_up = "low";

dffeas \dffe7a[3] (
	.clk(clock0),
	.d(\dffe7a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_3),
	.prn(vcc));
defparam \dffe7a[3] .is_wysiwyg = "true";
defparam \dffe7a[3] .power_up = "low";

dffeas \dffe7a[2] (
	.clk(clock0),
	.d(\dffe7a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_2),
	.prn(vcc));
defparam \dffe7a[2] .is_wysiwyg = "true";
defparam \dffe7a[2] .power_up = "low";

dffeas \dffe7a[1] (
	.clk(clock0),
	.d(\dffe7a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_1),
	.prn(vcc));
defparam \dffe7a[1] .is_wysiwyg = "true";
defparam \dffe7a[1] .power_up = "low";

dffeas \dffe7a[0] (
	.clk(clock0),
	.d(\dffe7a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_0),
	.prn(vcc));
defparam \dffe7a[0] .is_wysiwyg = "true";
defparam \dffe7a[0] .power_up = "low";

dffeas \dffe7a[19] (
	.clk(clock0),
	.d(\dffe7a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_19),
	.prn(vcc));
defparam \dffe7a[19] .is_wysiwyg = "true";
defparam \dffe7a[19] .power_up = "low";

dffeas \dffe7a[18] (
	.clk(clock0),
	.d(\dffe7a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_18),
	.prn(vcc));
defparam \dffe7a[18] .is_wysiwyg = "true";
defparam \dffe7a[18] .power_up = "low";

dffeas \dffe7a[17] (
	.clk(clock0),
	.d(\dffe7a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_17),
	.prn(vcc));
defparam \dffe7a[17] .is_wysiwyg = "true";
defparam \dffe7a[17] .power_up = "low";

dffeas \dffe7a[16] (
	.clk(clock0),
	.d(\dffe7a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_16),
	.prn(vcc));
defparam \dffe7a[16] .is_wysiwyg = "true";
defparam \dffe7a[16] .power_up = "low";

cycloneive_lcell_comb \dffe7a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe7a[0]~20_combout ),
	.cout(\dffe7a[0]~21 ));
defparam \dffe7a[0]~20 .lut_mask = 16'h66DD;
defparam \dffe7a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe7a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[0]~21 ),
	.combout(\dffe7a[1]~22_combout ),
	.cout(\dffe7a[1]~23 ));
defparam \dffe7a[1]~22 .lut_mask = 16'h96BF;
defparam \dffe7a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[1]~23 ),
	.combout(\dffe7a[2]~24_combout ),
	.cout(\dffe7a[2]~25 ));
defparam \dffe7a[2]~24 .lut_mask = 16'h96DF;
defparam \dffe7a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[2]~25 ),
	.combout(\dffe7a[3]~26_combout ),
	.cout(\dffe7a[3]~27 ));
defparam \dffe7a[3]~26 .lut_mask = 16'h96BF;
defparam \dffe7a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[3]~27 ),
	.combout(\dffe7a[4]~28_combout ),
	.cout(\dffe7a[4]~29 ));
defparam \dffe7a[4]~28 .lut_mask = 16'h96DF;
defparam \dffe7a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[4]~29 ),
	.combout(\dffe7a[5]~30_combout ),
	.cout(\dffe7a[5]~31 ));
defparam \dffe7a[5]~30 .lut_mask = 16'h96BF;
defparam \dffe7a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[5]~31 ),
	.combout(\dffe7a[6]~32_combout ),
	.cout(\dffe7a[6]~33 ));
defparam \dffe7a[6]~32 .lut_mask = 16'h96DF;
defparam \dffe7a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[6]~33 ),
	.combout(\dffe7a[7]~34_combout ),
	.cout(\dffe7a[7]~35 ));
defparam \dffe7a[7]~34 .lut_mask = 16'h96BF;
defparam \dffe7a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[7]~35 ),
	.combout(\dffe7a[8]~36_combout ),
	.cout(\dffe7a[8]~37 ));
defparam \dffe7a[8]~36 .lut_mask = 16'h96DF;
defparam \dffe7a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[8]~37 ),
	.combout(\dffe7a[9]~38_combout ),
	.cout(\dffe7a[9]~39 ));
defparam \dffe7a[9]~38 .lut_mask = 16'h96BF;
defparam \dffe7a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[9]~39 ),
	.combout(\dffe7a[10]~40_combout ),
	.cout(\dffe7a[10]~41 ));
defparam \dffe7a[10]~40 .lut_mask = 16'h96DF;
defparam \dffe7a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[10]~41 ),
	.combout(\dffe7a[11]~42_combout ),
	.cout(\dffe7a[11]~43 ));
defparam \dffe7a[11]~42 .lut_mask = 16'h96BF;
defparam \dffe7a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[11]~43 ),
	.combout(\dffe7a[12]~44_combout ),
	.cout(\dffe7a[12]~45 ));
defparam \dffe7a[12]~44 .lut_mask = 16'h96DF;
defparam \dffe7a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[12]~45 ),
	.combout(\dffe7a[13]~46_combout ),
	.cout(\dffe7a[13]~47 ));
defparam \dffe7a[13]~46 .lut_mask = 16'h96BF;
defparam \dffe7a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[13]~47 ),
	.combout(\dffe7a[14]~48_combout ),
	.cout(\dffe7a[14]~49 ));
defparam \dffe7a[14]~48 .lut_mask = 16'h96DF;
defparam \dffe7a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[14]~49 ),
	.combout(\dffe7a[15]~50_combout ),
	.cout(\dffe7a[15]~51 ));
defparam \dffe7a[15]~50 .lut_mask = 16'h96BF;
defparam \dffe7a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[15]~51 ),
	.combout(\dffe7a[16]~52_combout ),
	.cout(\dffe7a[16]~53 ));
defparam \dffe7a[16]~52 .lut_mask = 16'h96DF;
defparam \dffe7a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[16]~53 ),
	.combout(\dffe7a[17]~54_combout ),
	.cout(\dffe7a[17]~55 ));
defparam \dffe7a[17]~54 .lut_mask = 16'h96BF;
defparam \dffe7a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[17]~55 ),
	.combout(\dffe7a[18]~56_combout ),
	.cout(\dffe7a[18]~57 ));
defparam \dffe7a[18]~56 .lut_mask = 16'h96DF;
defparam \dffe7a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe7a[18]~57 ),
	.combout(\dffe7a[19]~58_combout ),
	.cout());
defparam \dffe7a[19]~58 .lut_mask = 16'h9696;
defparam \dffe7a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91_6 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_7 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_pround_2 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_3 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_3 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj_2 auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj_2 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_r_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_r_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_r_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_r_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_r_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_r_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_r_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_r_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_r_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_r_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_r_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_r_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_r_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_r_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_r_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_r_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_r_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_r_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_r_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_3 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_4 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_4 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj_3 auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj_3 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_i_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_i_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_i_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_i_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_i_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_i_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_i_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_i_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_i_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_i_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_i_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_i_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_i_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_i_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_i_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_i_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_i_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_i_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_i_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm2|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_tdl_2 (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_tdl_3 (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_cmult_std_2 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_5_11,
	tdl_arr_9_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_7_1,
	tdl_arr_7_11,
	tdl_arr_8_1,
	tdl_arr_8_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_3_1,
	tdl_arr_3_11,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk)/* synthesis synthesis_greybox=1 */;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_5_11;
output 	tdl_arr_9_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_7_1;
output 	tdl_arr_7_11;
output 	tdl_arr_8_1;
output 	tdl_arr_8_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_3_1;
output 	tdl_arr_3_11;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ;
wire \gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ;
wire \gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \result_i_tmp[15]~q ;
wire \result_i_tmp[14]~q ;
wire \result_i_tmp[13]~q ;
wire \result_i_tmp[12]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[10]~q ;
wire \result_i_tmp[9]~q ;
wire \result_i_tmp[8]~q ;
wire \result_i_tmp[7]~q ;
wire \result_i_tmp[6]~q ;
wire \result_i_tmp[5]~q ;
wire \result_i_tmp[4]~q ;
wire \result_i_tmp[3]~q ;
wire \result_i_tmp[2]~q ;
wire \result_i_tmp[1]~q ;
wire \result_i_tmp[0]~q ;
wire \result_i_tmp[19]~q ;
wire \result_i_tmp[18]~q ;
wire \result_i_tmp[17]~q ;
wire \result_i_tmp[16]~q ;
wire \result_r_tmp[15]~q ;
wire \result_r_tmp[14]~q ;
wire \result_r_tmp[13]~q ;
wire \result_r_tmp[12]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[10]~q ;
wire \result_r_tmp[9]~q ;
wire \result_r_tmp[8]~q ;
wire \result_r_tmp[7]~q ;
wire \result_r_tmp[6]~q ;
wire \result_r_tmp[5]~q ;
wire \result_r_tmp[4]~q ;
wire \result_r_tmp[3]~q ;
wire \result_r_tmp[2]~q ;
wire \result_r_tmp[1]~q ;
wire \result_r_tmp[0]~q ;
wire \result_r_tmp[19]~q ;
wire \result_r_tmp[18]~q ;
wire \result_r_tmp[17]~q ;
wire \result_r_tmp[16]~q ;


fftsign_asj_fft_tdl_4 \gen_ma:gen_ma_full:imag_delay (
	.data_in({\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_9_1(tdl_arr_9_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_8_1(tdl_arr_8_1),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_3_1(tdl_arr_3_1),
	.clk(clk));

fftsign_asj_fft_tdl_5 \gen_ma:gen_ma_full:real_delay (
	.data_in({\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,
\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q }),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_9_1(tdl_arr_9_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_8_1(tdl_arr_8_11),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_3_1(tdl_arr_3_11),
	.clk(clk));

fftsign_asj_fft_pround_5 \gen_ma:gen_ma_full:u1 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.result_i_tmp_19(\result_i_tmp[19]~q ),
	.result_i_tmp_18(\result_i_tmp[18]~q ),
	.result_i_tmp_17(\result_i_tmp[17]~q ),
	.result_i_tmp_16(\result_i_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_pround_4 \gen_ma:gen_ma_full:u0 (
	.pipeline_dffe_15(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_19(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_16(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_12(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_14(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.global_clock_enable(global_clock_enable),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.result_r_tmp_19(\result_r_tmp[19]~q ),
	.result_r_tmp_18(\result_r_tmp[18]~q ),
	.result_r_tmp_17(\result_r_tmp[17]~q ),
	.result_r_tmp_16(\result_r_tmp[16]~q ),
	.clk(clk));

fftsign_asj_fft_mult_add_4 \gen_ma:gen_ma_full:ma (
	.dffe5a_15(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.dffe5a_14(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.dffe5a_13(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.dffe5a_12(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.dffe5a_11(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.dffe5a_10(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.dffe5a_9(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.dffe5a_8(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.dffe5a_7(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.dffe5a_6(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.dffe5a_5(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.dffe5a_4(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.dffe5a_3(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.dffe5a_2(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.dffe5a_1(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.dffe5a_0(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.dffe5a_19(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.dffe5a_18(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.dffe5a_17(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.dffe5a_16(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.twiddle_data218(twiddle_data218),
	.twiddle_data219(twiddle_data219),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data208(twiddle_data208),
	.twiddle_data209(twiddle_data209),
	.clk(clk));

fftsign_asj_fft_mult_add_5 \gen_ma:gen_ma_full:ms (
	.dffe7a_15(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.dffe7a_14(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.dffe7a_13(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.dffe7a_12(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.dffe7a_11(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.dffe7a_10(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.dffe7a_9(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.dffe7a_8(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.dffe7a_7(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.dffe7a_6(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.dffe7a_5(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.dffe7a_4(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.dffe7a_3(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.dffe7a_2(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.dffe7a_1(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.dffe7a_0(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.dffe7a_19(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.dffe7a_18(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.dffe7a_17(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.dffe7a_16(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.twiddle_data218(twiddle_data218),
	.twiddle_data219(twiddle_data219),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data208(twiddle_data208),
	.twiddle_data209(twiddle_data209),
	.clk(clk));

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

dffeas \result_i_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[19]~q ),
	.prn(vcc));
defparam \result_i_tmp[19] .is_wysiwyg = "true";
defparam \result_i_tmp[19] .power_up = "low";

dffeas \result_i_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[18]~q ),
	.prn(vcc));
defparam \result_i_tmp[18] .is_wysiwyg = "true";
defparam \result_i_tmp[18] .power_up = "low";

dffeas \result_i_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[17]~q ),
	.prn(vcc));
defparam \result_i_tmp[17] .is_wysiwyg = "true";
defparam \result_i_tmp[17] .power_up = "low";

dffeas \result_i_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ma|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_i_tmp[16]~q ),
	.prn(vcc));
defparam \result_i_tmp[16] .is_wysiwyg = "true";
defparam \result_i_tmp[16] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

dffeas \result_r_tmp[19] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[19]~q ),
	.prn(vcc));
defparam \result_r_tmp[19] .is_wysiwyg = "true";
defparam \result_r_tmp[19] .power_up = "low";

dffeas \result_r_tmp[18] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[18]~q ),
	.prn(vcc));
defparam \result_r_tmp[18] .is_wysiwyg = "true";
defparam \result_r_tmp[18] .power_up = "low";

dffeas \result_r_tmp[17] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[17]~q ),
	.prn(vcc));
defparam \result_r_tmp[17] .is_wysiwyg = "true";
defparam \result_r_tmp[17] .power_up = "low";

dffeas \result_r_tmp[16] (
	.clk(clk),
	.d(\gen_ma:gen_ma_full:ms|MULT_ADD_component|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_r_tmp[16]~q ),
	.prn(vcc));
defparam \result_r_tmp[16] .is_wysiwyg = "true";
defparam \result_r_tmp[16] .power_up = "low";

endmodule

module fftsign_asj_fft_mult_add_4 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_4 MULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.twiddle_data218(twiddle_data218),
	.twiddle_data219(twiddle_data219),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data208(twiddle_data208),
	.twiddle_data209(twiddle_data209),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add_4 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old_4 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2,pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,
pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.ena0(global_clock_enable),
	.datab({twiddle_data219,twiddle_data218,twiddle_data217,twiddle_data216,twiddle_data215,twiddle_data214,twiddle_data213,twiddle_data212,twiddle_data211,twiddle_data210,twiddle_data209,twiddle_data208,twiddle_data207,twiddle_data206,twiddle_data205,twiddle_data204,twiddle_data203,
twiddle_data202,twiddle_data201,twiddle_data200}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old_4 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_5 ALTMULT_ADD_component(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_5 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_kk6g_2 auto_generated(
	.dffe5a_15(dffe5a_15),
	.dffe5a_14(dffe5a_14),
	.dffe5a_13(dffe5a_13),
	.dffe5a_12(dffe5a_12),
	.dffe5a_11(dffe5a_11),
	.dffe5a_10(dffe5a_10),
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_5(dffe5a_5),
	.dffe5a_4(dffe5a_4),
	.dffe5a_3(dffe5a_3),
	.dffe5a_2(dffe5a_2),
	.dffe5a_1(dffe5a_1),
	.dffe5a_0(dffe5a_0),
	.dffe5a_19(dffe5a_19),
	.dffe5a_18(dffe5a_18),
	.dffe5a_17(dffe5a_17),
	.dffe5a_16(dffe5a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_kk6g_2 (
	dffe5a_15,
	dffe5a_14,
	dffe5a_13,
	dffe5a_12,
	dffe5a_11,
	dffe5a_10,
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_5,
	dffe5a_4,
	dffe5a_3,
	dffe5a_2,
	dffe5a_1,
	dffe5a_0,
	dffe5a_19,
	dffe5a_18,
	dffe5a_17,
	dffe5a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_15;
output 	dffe5a_14;
output 	dffe5a_13;
output 	dffe5a_12;
output 	dffe5a_11;
output 	dffe5a_10;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_5;
output 	dffe5a_4;
output 	dffe5a_3;
output 	dffe5a_2;
output 	dffe5a_1;
output 	dffe5a_0;
output 	dffe5a_19;
output 	dffe5a_18;
output 	dffe5a_17;
output 	dffe5a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe5a[0]~21 ;
wire \dffe5a[1]~23 ;
wire \dffe5a[2]~25 ;
wire \dffe5a[3]~27 ;
wire \dffe5a[4]~29 ;
wire \dffe5a[5]~31 ;
wire \dffe5a[6]~33 ;
wire \dffe5a[7]~35 ;
wire \dffe5a[8]~37 ;
wire \dffe5a[9]~39 ;
wire \dffe5a[10]~41 ;
wire \dffe5a[11]~43 ;
wire \dffe5a[12]~45 ;
wire \dffe5a[13]~47 ;
wire \dffe5a[14]~49 ;
wire \dffe5a[15]~50_combout ;
wire \dffe5a[14]~48_combout ;
wire \dffe5a[13]~46_combout ;
wire \dffe5a[12]~44_combout ;
wire \dffe5a[11]~42_combout ;
wire \dffe5a[10]~40_combout ;
wire \dffe5a[9]~38_combout ;
wire \dffe5a[8]~36_combout ;
wire \dffe5a[7]~34_combout ;
wire \dffe5a[6]~32_combout ;
wire \dffe5a[5]~30_combout ;
wire \dffe5a[4]~28_combout ;
wire \dffe5a[3]~26_combout ;
wire \dffe5a[2]~24_combout ;
wire \dffe5a[1]~22_combout ;
wire \dffe5a[0]~20_combout ;
wire \dffe5a[15]~51 ;
wire \dffe5a[16]~53 ;
wire \dffe5a[17]~55 ;
wire \dffe5a[18]~57 ;
wire \dffe5a[19]~58_combout ;
wire \dffe5a[18]~56_combout ;
wire \dffe5a[17]~54_combout ;
wire \dffe5a[16]~52_combout ;


fftsign_ded_mult_9a91_9 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91_8 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe5a[15] (
	.clk(clock0),
	.d(\dffe5a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_15),
	.prn(vcc));
defparam \dffe5a[15] .is_wysiwyg = "true";
defparam \dffe5a[15] .power_up = "low";

dffeas \dffe5a[14] (
	.clk(clock0),
	.d(\dffe5a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_14),
	.prn(vcc));
defparam \dffe5a[14] .is_wysiwyg = "true";
defparam \dffe5a[14] .power_up = "low";

dffeas \dffe5a[13] (
	.clk(clock0),
	.d(\dffe5a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_13),
	.prn(vcc));
defparam \dffe5a[13] .is_wysiwyg = "true";
defparam \dffe5a[13] .power_up = "low";

dffeas \dffe5a[12] (
	.clk(clock0),
	.d(\dffe5a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_12),
	.prn(vcc));
defparam \dffe5a[12] .is_wysiwyg = "true";
defparam \dffe5a[12] .power_up = "low";

dffeas \dffe5a[11] (
	.clk(clock0),
	.d(\dffe5a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_11),
	.prn(vcc));
defparam \dffe5a[11] .is_wysiwyg = "true";
defparam \dffe5a[11] .power_up = "low";

dffeas \dffe5a[10] (
	.clk(clock0),
	.d(\dffe5a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_10),
	.prn(vcc));
defparam \dffe5a[10] .is_wysiwyg = "true";
defparam \dffe5a[10] .power_up = "low";

dffeas \dffe5a[9] (
	.clk(clock0),
	.d(\dffe5a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_9),
	.prn(vcc));
defparam \dffe5a[9] .is_wysiwyg = "true";
defparam \dffe5a[9] .power_up = "low";

dffeas \dffe5a[8] (
	.clk(clock0),
	.d(\dffe5a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_8),
	.prn(vcc));
defparam \dffe5a[8] .is_wysiwyg = "true";
defparam \dffe5a[8] .power_up = "low";

dffeas \dffe5a[7] (
	.clk(clock0),
	.d(\dffe5a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_7),
	.prn(vcc));
defparam \dffe5a[7] .is_wysiwyg = "true";
defparam \dffe5a[7] .power_up = "low";

dffeas \dffe5a[6] (
	.clk(clock0),
	.d(\dffe5a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_6),
	.prn(vcc));
defparam \dffe5a[6] .is_wysiwyg = "true";
defparam \dffe5a[6] .power_up = "low";

dffeas \dffe5a[5] (
	.clk(clock0),
	.d(\dffe5a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_5),
	.prn(vcc));
defparam \dffe5a[5] .is_wysiwyg = "true";
defparam \dffe5a[5] .power_up = "low";

dffeas \dffe5a[4] (
	.clk(clock0),
	.d(\dffe5a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_4),
	.prn(vcc));
defparam \dffe5a[4] .is_wysiwyg = "true";
defparam \dffe5a[4] .power_up = "low";

dffeas \dffe5a[3] (
	.clk(clock0),
	.d(\dffe5a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_3),
	.prn(vcc));
defparam \dffe5a[3] .is_wysiwyg = "true";
defparam \dffe5a[3] .power_up = "low";

dffeas \dffe5a[2] (
	.clk(clock0),
	.d(\dffe5a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_2),
	.prn(vcc));
defparam \dffe5a[2] .is_wysiwyg = "true";
defparam \dffe5a[2] .power_up = "low";

dffeas \dffe5a[1] (
	.clk(clock0),
	.d(\dffe5a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_1),
	.prn(vcc));
defparam \dffe5a[1] .is_wysiwyg = "true";
defparam \dffe5a[1] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock0),
	.d(\dffe5a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_0),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

dffeas \dffe5a[19] (
	.clk(clock0),
	.d(\dffe5a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_19),
	.prn(vcc));
defparam \dffe5a[19] .is_wysiwyg = "true";
defparam \dffe5a[19] .power_up = "low";

dffeas \dffe5a[18] (
	.clk(clock0),
	.d(\dffe5a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_18),
	.prn(vcc));
defparam \dffe5a[18] .is_wysiwyg = "true";
defparam \dffe5a[18] .power_up = "low";

dffeas \dffe5a[17] (
	.clk(clock0),
	.d(\dffe5a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_17),
	.prn(vcc));
defparam \dffe5a[17] .is_wysiwyg = "true";
defparam \dffe5a[17] .power_up = "low";

dffeas \dffe5a[16] (
	.clk(clock0),
	.d(\dffe5a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_16),
	.prn(vcc));
defparam \dffe5a[16] .is_wysiwyg = "true";
defparam \dffe5a[16] .power_up = "low";

cycloneive_lcell_comb \dffe5a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe5a[0]~20_combout ),
	.cout(\dffe5a[0]~21 ));
defparam \dffe5a[0]~20 .lut_mask = 16'h66EE;
defparam \dffe5a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe5a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[0]~21 ),
	.combout(\dffe5a[1]~22_combout ),
	.cout(\dffe5a[1]~23 ));
defparam \dffe5a[1]~22 .lut_mask = 16'h967F;
defparam \dffe5a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[1]~23 ),
	.combout(\dffe5a[2]~24_combout ),
	.cout(\dffe5a[2]~25 ));
defparam \dffe5a[2]~24 .lut_mask = 16'h96EF;
defparam \dffe5a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[2]~25 ),
	.combout(\dffe5a[3]~26_combout ),
	.cout(\dffe5a[3]~27 ));
defparam \dffe5a[3]~26 .lut_mask = 16'h967F;
defparam \dffe5a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[3]~27 ),
	.combout(\dffe5a[4]~28_combout ),
	.cout(\dffe5a[4]~29 ));
defparam \dffe5a[4]~28 .lut_mask = 16'h96EF;
defparam \dffe5a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[4]~29 ),
	.combout(\dffe5a[5]~30_combout ),
	.cout(\dffe5a[5]~31 ));
defparam \dffe5a[5]~30 .lut_mask = 16'h967F;
defparam \dffe5a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[5]~31 ),
	.combout(\dffe5a[6]~32_combout ),
	.cout(\dffe5a[6]~33 ));
defparam \dffe5a[6]~32 .lut_mask = 16'h96EF;
defparam \dffe5a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[6]~33 ),
	.combout(\dffe5a[7]~34_combout ),
	.cout(\dffe5a[7]~35 ));
defparam \dffe5a[7]~34 .lut_mask = 16'h967F;
defparam \dffe5a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[7]~35 ),
	.combout(\dffe5a[8]~36_combout ),
	.cout(\dffe5a[8]~37 ));
defparam \dffe5a[8]~36 .lut_mask = 16'h96EF;
defparam \dffe5a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[8]~37 ),
	.combout(\dffe5a[9]~38_combout ),
	.cout(\dffe5a[9]~39 ));
defparam \dffe5a[9]~38 .lut_mask = 16'h967F;
defparam \dffe5a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[9]~39 ),
	.combout(\dffe5a[10]~40_combout ),
	.cout(\dffe5a[10]~41 ));
defparam \dffe5a[10]~40 .lut_mask = 16'h96EF;
defparam \dffe5a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[10]~41 ),
	.combout(\dffe5a[11]~42_combout ),
	.cout(\dffe5a[11]~43 ));
defparam \dffe5a[11]~42 .lut_mask = 16'h967F;
defparam \dffe5a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[11]~43 ),
	.combout(\dffe5a[12]~44_combout ),
	.cout(\dffe5a[12]~45 ));
defparam \dffe5a[12]~44 .lut_mask = 16'h96EF;
defparam \dffe5a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[12]~45 ),
	.combout(\dffe5a[13]~46_combout ),
	.cout(\dffe5a[13]~47 ));
defparam \dffe5a[13]~46 .lut_mask = 16'h967F;
defparam \dffe5a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[13]~47 ),
	.combout(\dffe5a[14]~48_combout ),
	.cout(\dffe5a[14]~49 ));
defparam \dffe5a[14]~48 .lut_mask = 16'h96EF;
defparam \dffe5a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[14]~49 ),
	.combout(\dffe5a[15]~50_combout ),
	.cout(\dffe5a[15]~51 ));
defparam \dffe5a[15]~50 .lut_mask = 16'h967F;
defparam \dffe5a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[15]~51 ),
	.combout(\dffe5a[16]~52_combout ),
	.cout(\dffe5a[16]~53 ));
defparam \dffe5a[16]~52 .lut_mask = 16'h96EF;
defparam \dffe5a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[16]~53 ),
	.combout(\dffe5a[17]~54_combout ),
	.cout(\dffe5a[17]~55 ));
defparam \dffe5a[17]~54 .lut_mask = 16'h967F;
defparam \dffe5a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[17]~55 ),
	.combout(\dffe5a[18]~56_combout ),
	.cout(\dffe5a[18]~57 ));
defparam \dffe5a[18]~56 .lut_mask = 16'h96EF;
defparam \dffe5a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe5a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe5a[18]~57 ),
	.combout(\dffe5a[19]~58_combout ),
	.cout());
defparam \dffe5a[19]~58 .lut_mask = 16'h9696;
defparam \dffe5a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91_8 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_9 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_mult_add_5 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_5 MULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_41(pipeline_dffe_41),
	.pipeline_dffe_51(pipeline_dffe_51),
	.pipeline_dffe_61(pipeline_dffe_61),
	.pipeline_dffe_71(pipeline_dffe_71),
	.pipeline_dffe_81(pipeline_dffe_81),
	.pipeline_dffe_91(pipeline_dffe_91),
	.pipeline_dffe_101(pipeline_dffe_101),
	.pipeline_dffe_111(pipeline_dffe_111),
	.global_clock_enable(global_clock_enable),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.twiddle_data218(twiddle_data218),
	.twiddle_data219(twiddle_data219),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.twiddle_data207(twiddle_data207),
	.twiddle_data208(twiddle_data208),
	.twiddle_data209(twiddle_data209),
	.clk(clk));

endmodule

module fftsign_altera_fft_mult_add_5 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	global_clock_enable,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	twiddle_data218,
	twiddle_data219,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	twiddle_data207,
	twiddle_data208,
	twiddle_data209,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	global_clock_enable;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	twiddle_data218;
input 	twiddle_data219;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	twiddle_data207;
input 	twiddle_data208;
input 	twiddle_data209;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altera_fft_mult_add_old_5 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({pipeline_dffe_111,pipeline_dffe_101,pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21,pipeline_dffe_11,pipeline_dffe_10,pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,
pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.ena0(global_clock_enable),
	.datab({twiddle_data219,twiddle_data218,twiddle_data217,twiddle_data216,twiddle_data215,twiddle_data214,twiddle_data213,twiddle_data212,twiddle_data211,twiddle_data210,twiddle_data209,twiddle_data208,twiddle_data207,twiddle_data206,twiddle_data205,twiddle_data204,twiddle_data203,
twiddle_data202,twiddle_data201,twiddle_data200}),
	.clock0(clk));

endmodule

module fftsign_altera_fft_mult_add_old_5 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_altmult_add_6 ALTMULT_ADD_component(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_altmult_add_6 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_mult_add_ll6g_2 auto_generated(
	.dffe7a_15(dffe7a_15),
	.dffe7a_14(dffe7a_14),
	.dffe7a_13(dffe7a_13),
	.dffe7a_12(dffe7a_12),
	.dffe7a_11(dffe7a_11),
	.dffe7a_10(dffe7a_10),
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_5(dffe7a_5),
	.dffe7a_4(dffe7a_4),
	.dffe7a_3(dffe7a_3),
	.dffe7a_2(dffe7a_2),
	.dffe7a_1(dffe7a_1),
	.dffe7a_0(dffe7a_0),
	.dffe7a_19(dffe7a_19),
	.dffe7a_18(dffe7a_18),
	.dffe7a_17(dffe7a_17),
	.dffe7a_16(dffe7a_16),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena0(ena0),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock0(clock0));

endmodule

module fftsign_mult_add_ll6g_2 (
	dffe7a_15,
	dffe7a_14,
	dffe7a_13,
	dffe7a_12,
	dffe7a_11,
	dffe7a_10,
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_5,
	dffe7a_4,
	dffe7a_3,
	dffe7a_2,
	dffe7a_1,
	dffe7a_0,
	dffe7a_19,
	dffe7a_18,
	dffe7a_17,
	dffe7a_16,
	dataa,
	ena0,
	datab,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_15;
output 	dffe7a_14;
output 	dffe7a_13;
output 	dffe7a_12;
output 	dffe7a_11;
output 	dffe7a_10;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_5;
output 	dffe7a_4;
output 	dffe7a_3;
output 	dffe7a_2;
output 	dffe7a_1;
output 	dffe7a_0;
output 	dffe7a_19;
output 	dffe7a_18;
output 	dffe7a_17;
output 	dffe7a_16;
input 	[19:0] dataa;
input 	ena0;
input 	[19:0] datab;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult2|mac_out9~DATAOUT16 ;
wire \ded_mult2|mac_out9~DATAOUT17 ;
wire \ded_mult2|mac_out9~DATAOUT18 ;
wire \ded_mult2|mac_out9~DATAOUT19 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~DATAOUT16 ;
wire \ded_mult1|mac_out9~DATAOUT17 ;
wire \ded_mult1|mac_out9~DATAOUT18 ;
wire \ded_mult1|mac_out9~DATAOUT19 ;
wire \dffe7a[0]~21 ;
wire \dffe7a[1]~23 ;
wire \dffe7a[2]~25 ;
wire \dffe7a[3]~27 ;
wire \dffe7a[4]~29 ;
wire \dffe7a[5]~31 ;
wire \dffe7a[6]~33 ;
wire \dffe7a[7]~35 ;
wire \dffe7a[8]~37 ;
wire \dffe7a[9]~39 ;
wire \dffe7a[10]~41 ;
wire \dffe7a[11]~43 ;
wire \dffe7a[12]~45 ;
wire \dffe7a[13]~47 ;
wire \dffe7a[14]~49 ;
wire \dffe7a[15]~50_combout ;
wire \dffe7a[14]~48_combout ;
wire \dffe7a[13]~46_combout ;
wire \dffe7a[12]~44_combout ;
wire \dffe7a[11]~42_combout ;
wire \dffe7a[10]~40_combout ;
wire \dffe7a[9]~38_combout ;
wire \dffe7a[8]~36_combout ;
wire \dffe7a[7]~34_combout ;
wire \dffe7a[6]~32_combout ;
wire \dffe7a[5]~30_combout ;
wire \dffe7a[4]~28_combout ;
wire \dffe7a[3]~26_combout ;
wire \dffe7a[2]~24_combout ;
wire \dffe7a[1]~22_combout ;
wire \dffe7a[0]~20_combout ;
wire \dffe7a[15]~51 ;
wire \dffe7a[16]~53 ;
wire \dffe7a[17]~55 ;
wire \dffe7a[18]~57 ;
wire \dffe7a[19]~58_combout ;
wire \dffe7a[18]~56_combout ;
wire \dffe7a[17]~54_combout ;
wire \dffe7a[16]~52_combout ;


fftsign_ded_mult_9a91_11 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult2|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult2|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult2|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult2|mac_out9~DATAOUT19 ),
	.dataa({dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10]}),
	.clock({gnd,gnd,gnd,clock0}));

fftsign_ded_mult_9a91_10 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.mac_out917(\ded_mult1|mac_out9~DATAOUT16 ),
	.mac_out918(\ded_mult1|mac_out9~DATAOUT17 ),
	.mac_out919(\ded_mult1|mac_out9~DATAOUT18 ),
	.mac_out920(\ded_mult1|mac_out9~DATAOUT19 ),
	.dataa({dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.clock({gnd,gnd,gnd,clock0}));

dffeas \dffe7a[15] (
	.clk(clock0),
	.d(\dffe7a[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_15),
	.prn(vcc));
defparam \dffe7a[15] .is_wysiwyg = "true";
defparam \dffe7a[15] .power_up = "low";

dffeas \dffe7a[14] (
	.clk(clock0),
	.d(\dffe7a[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_14),
	.prn(vcc));
defparam \dffe7a[14] .is_wysiwyg = "true";
defparam \dffe7a[14] .power_up = "low";

dffeas \dffe7a[13] (
	.clk(clock0),
	.d(\dffe7a[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_13),
	.prn(vcc));
defparam \dffe7a[13] .is_wysiwyg = "true";
defparam \dffe7a[13] .power_up = "low";

dffeas \dffe7a[12] (
	.clk(clock0),
	.d(\dffe7a[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_12),
	.prn(vcc));
defparam \dffe7a[12] .is_wysiwyg = "true";
defparam \dffe7a[12] .power_up = "low";

dffeas \dffe7a[11] (
	.clk(clock0),
	.d(\dffe7a[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_11),
	.prn(vcc));
defparam \dffe7a[11] .is_wysiwyg = "true";
defparam \dffe7a[11] .power_up = "low";

dffeas \dffe7a[10] (
	.clk(clock0),
	.d(\dffe7a[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_10),
	.prn(vcc));
defparam \dffe7a[10] .is_wysiwyg = "true";
defparam \dffe7a[10] .power_up = "low";

dffeas \dffe7a[9] (
	.clk(clock0),
	.d(\dffe7a[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_9),
	.prn(vcc));
defparam \dffe7a[9] .is_wysiwyg = "true";
defparam \dffe7a[9] .power_up = "low";

dffeas \dffe7a[8] (
	.clk(clock0),
	.d(\dffe7a[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_8),
	.prn(vcc));
defparam \dffe7a[8] .is_wysiwyg = "true";
defparam \dffe7a[8] .power_up = "low";

dffeas \dffe7a[7] (
	.clk(clock0),
	.d(\dffe7a[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_7),
	.prn(vcc));
defparam \dffe7a[7] .is_wysiwyg = "true";
defparam \dffe7a[7] .power_up = "low";

dffeas \dffe7a[6] (
	.clk(clock0),
	.d(\dffe7a[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_6),
	.prn(vcc));
defparam \dffe7a[6] .is_wysiwyg = "true";
defparam \dffe7a[6] .power_up = "low";

dffeas \dffe7a[5] (
	.clk(clock0),
	.d(\dffe7a[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_5),
	.prn(vcc));
defparam \dffe7a[5] .is_wysiwyg = "true";
defparam \dffe7a[5] .power_up = "low";

dffeas \dffe7a[4] (
	.clk(clock0),
	.d(\dffe7a[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_4),
	.prn(vcc));
defparam \dffe7a[4] .is_wysiwyg = "true";
defparam \dffe7a[4] .power_up = "low";

dffeas \dffe7a[3] (
	.clk(clock0),
	.d(\dffe7a[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_3),
	.prn(vcc));
defparam \dffe7a[3] .is_wysiwyg = "true";
defparam \dffe7a[3] .power_up = "low";

dffeas \dffe7a[2] (
	.clk(clock0),
	.d(\dffe7a[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_2),
	.prn(vcc));
defparam \dffe7a[2] .is_wysiwyg = "true";
defparam \dffe7a[2] .power_up = "low";

dffeas \dffe7a[1] (
	.clk(clock0),
	.d(\dffe7a[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_1),
	.prn(vcc));
defparam \dffe7a[1] .is_wysiwyg = "true";
defparam \dffe7a[1] .power_up = "low";

dffeas \dffe7a[0] (
	.clk(clock0),
	.d(\dffe7a[0]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_0),
	.prn(vcc));
defparam \dffe7a[0] .is_wysiwyg = "true";
defparam \dffe7a[0] .power_up = "low";

dffeas \dffe7a[19] (
	.clk(clock0),
	.d(\dffe7a[19]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_19),
	.prn(vcc));
defparam \dffe7a[19] .is_wysiwyg = "true";
defparam \dffe7a[19] .power_up = "low";

dffeas \dffe7a[18] (
	.clk(clock0),
	.d(\dffe7a[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_18),
	.prn(vcc));
defparam \dffe7a[18] .is_wysiwyg = "true";
defparam \dffe7a[18] .power_up = "low";

dffeas \dffe7a[17] (
	.clk(clock0),
	.d(\dffe7a[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_17),
	.prn(vcc));
defparam \dffe7a[17] .is_wysiwyg = "true";
defparam \dffe7a[17] .power_up = "low";

dffeas \dffe7a[16] (
	.clk(clock0),
	.d(\dffe7a[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_16),
	.prn(vcc));
defparam \dffe7a[16] .is_wysiwyg = "true";
defparam \dffe7a[16] .power_up = "low";

cycloneive_lcell_comb \dffe7a[0]~20 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe7a[0]~20_combout ),
	.cout(\dffe7a[0]~21 ));
defparam \dffe7a[0]~20 .lut_mask = 16'h66DD;
defparam \dffe7a[0]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe7a[1]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[0]~21 ),
	.combout(\dffe7a[1]~22_combout ),
	.cout(\dffe7a[1]~23 ));
defparam \dffe7a[1]~22 .lut_mask = 16'h96BF;
defparam \dffe7a[1]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[2]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[1]~23 ),
	.combout(\dffe7a[2]~24_combout ),
	.cout(\dffe7a[2]~25 ));
defparam \dffe7a[2]~24 .lut_mask = 16'h96DF;
defparam \dffe7a[2]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[3]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[2]~25 ),
	.combout(\dffe7a[3]~26_combout ),
	.cout(\dffe7a[3]~27 ));
defparam \dffe7a[3]~26 .lut_mask = 16'h96BF;
defparam \dffe7a[3]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[4]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[3]~27 ),
	.combout(\dffe7a[4]~28_combout ),
	.cout(\dffe7a[4]~29 ));
defparam \dffe7a[4]~28 .lut_mask = 16'h96DF;
defparam \dffe7a[4]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[5]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[4]~29 ),
	.combout(\dffe7a[5]~30_combout ),
	.cout(\dffe7a[5]~31 ));
defparam \dffe7a[5]~30 .lut_mask = 16'h96BF;
defparam \dffe7a[5]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[6]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[5]~31 ),
	.combout(\dffe7a[6]~32_combout ),
	.cout(\dffe7a[6]~33 ));
defparam \dffe7a[6]~32 .lut_mask = 16'h96DF;
defparam \dffe7a[6]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[7]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[6]~33 ),
	.combout(\dffe7a[7]~34_combout ),
	.cout(\dffe7a[7]~35 ));
defparam \dffe7a[7]~34 .lut_mask = 16'h96BF;
defparam \dffe7a[7]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[8]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[7]~35 ),
	.combout(\dffe7a[8]~36_combout ),
	.cout(\dffe7a[8]~37 ));
defparam \dffe7a[8]~36 .lut_mask = 16'h96DF;
defparam \dffe7a[8]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[9]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[8]~37 ),
	.combout(\dffe7a[9]~38_combout ),
	.cout(\dffe7a[9]~39 ));
defparam \dffe7a[9]~38 .lut_mask = 16'h96BF;
defparam \dffe7a[9]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[10]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[9]~39 ),
	.combout(\dffe7a[10]~40_combout ),
	.cout(\dffe7a[10]~41 ));
defparam \dffe7a[10]~40 .lut_mask = 16'h96DF;
defparam \dffe7a[10]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[11]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[10]~41 ),
	.combout(\dffe7a[11]~42_combout ),
	.cout(\dffe7a[11]~43 ));
defparam \dffe7a[11]~42 .lut_mask = 16'h96BF;
defparam \dffe7a[11]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[12]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[11]~43 ),
	.combout(\dffe7a[12]~44_combout ),
	.cout(\dffe7a[12]~45 ));
defparam \dffe7a[12]~44 .lut_mask = 16'h96DF;
defparam \dffe7a[12]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[13]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[12]~45 ),
	.combout(\dffe7a[13]~46_combout ),
	.cout(\dffe7a[13]~47 ));
defparam \dffe7a[13]~46 .lut_mask = 16'h96BF;
defparam \dffe7a[13]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[14]~48 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[13]~47 ),
	.combout(\dffe7a[14]~48_combout ),
	.cout(\dffe7a[14]~49 ));
defparam \dffe7a[14]~48 .lut_mask = 16'h96DF;
defparam \dffe7a[14]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[15]~50 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[14]~49 ),
	.combout(\dffe7a[15]~50_combout ),
	.cout(\dffe7a[15]~51 ));
defparam \dffe7a[15]~50 .lut_mask = 16'h96BF;
defparam \dffe7a[15]~50 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[16]~52 (
	.dataa(\ded_mult2|mac_out9~DATAOUT16 ),
	.datab(\ded_mult1|mac_out9~DATAOUT16 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[15]~51 ),
	.combout(\dffe7a[16]~52_combout ),
	.cout(\dffe7a[16]~53 ));
defparam \dffe7a[16]~52 .lut_mask = 16'h96DF;
defparam \dffe7a[16]~52 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[17]~54 (
	.dataa(\ded_mult2|mac_out9~DATAOUT17 ),
	.datab(\ded_mult1|mac_out9~DATAOUT17 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[16]~53 ),
	.combout(\dffe7a[17]~54_combout ),
	.cout(\dffe7a[17]~55 ));
defparam \dffe7a[17]~54 .lut_mask = 16'h96BF;
defparam \dffe7a[17]~54 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[18]~56 (
	.dataa(\ded_mult2|mac_out9~DATAOUT18 ),
	.datab(\ded_mult1|mac_out9~DATAOUT18 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[17]~55 ),
	.combout(\dffe7a[18]~56_combout ),
	.cout(\dffe7a[18]~57 ));
defparam \dffe7a[18]~56 .lut_mask = 16'h96DF;
defparam \dffe7a[18]~56 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dffe7a[19]~58 (
	.dataa(\ded_mult2|mac_out9~DATAOUT19 ),
	.datab(\ded_mult1|mac_out9~DATAOUT19 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe7a[18]~57 ),
	.combout(\dffe7a[19]~58_combout ),
	.cout());
defparam \dffe7a[19]~58 .lut_mask = 16'h9696;
defparam \dffe7a[19]~58 .sum_lutc_input = "cin";

endmodule

module fftsign_ded_mult_9a91_10 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_ded_mult_9a91_11 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	mac_out917,
	mac_out918,
	mac_out919,
	mac_out920,
	dataa,
	ena,
	datab,
	clock)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
output 	mac_out917;
output 	mac_out918;
output 	mac_out919;
output 	mac_out920;
input 	[9:0] dataa;
input 	[3:0] ena;
input 	[9:0] datab;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;
wire \mac_mult8~DATAOUT16 ;
wire \mac_mult8~DATAOUT17 ;
wire \mac_mult8~DATAOUT18 ;
wire \mac_mult8~DATAOUT19 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];
assign mac_out917 = mac_out9_DATAOUT_bus[16];
assign mac_out918 = mac_out9_DATAOUT_bus[17];
assign mac_out919 = mac_out9_DATAOUT_bus[18];
assign mac_out920 = mac_out9_DATAOUT_bus[19];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];
assign \mac_mult8~DATAOUT16  = mac_mult8_DATAOUT_bus[16];
assign \mac_mult8~DATAOUT17  = mac_mult8_DATAOUT_bus[17];
assign \mac_mult8~DATAOUT18  = mac_mult8_DATAOUT_bus[18];
assign \mac_mult8~DATAOUT19  = mac_mult8_DATAOUT_bus[19];

cycloneive_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT19 ,\mac_mult8~DATAOUT18 ,\mac_mult8~DATAOUT17 ,\mac_mult8~DATAOUT16 ,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,
\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 20;
defparam mac_out9.output_clock = "0";

cycloneive_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(gnd),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 10;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 10;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module fftsign_asj_fft_pround_4 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_5 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_5 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj_4 auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.result_r_tmp_8(result_r_tmp_8),
	.result_r_tmp_7(result_r_tmp_7),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.result_r_tmp_19(result_r_tmp_19),
	.result_r_tmp_18(result_r_tmp_18),
	.result_r_tmp_17(result_r_tmp_17),
	.result_r_tmp_16(result_r_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj_4 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_r_tmp_15,
	result_r_tmp_14,
	result_r_tmp_13,
	result_r_tmp_12,
	result_r_tmp_11,
	result_r_tmp_10,
	result_r_tmp_9,
	result_r_tmp_8,
	result_r_tmp_7,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	result_r_tmp_19,
	result_r_tmp_18,
	result_r_tmp_17,
	result_r_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_r_tmp_15;
input 	result_r_tmp_14;
input 	result_r_tmp_13;
input 	result_r_tmp_12;
input 	result_r_tmp_11;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
input 	result_r_tmp_8;
input 	result_r_tmp_7;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	result_r_tmp_19;
input 	result_r_tmp_18;
input 	result_r_tmp_17;
input 	result_r_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_r_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_r_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_r_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_r_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_r_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_r_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_r_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_r_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_r_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_r_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_r_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_r_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_r_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_r_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_r_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_r_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_r_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_r_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_r_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_r_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_5 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	global_clock_enable,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	global_clock_enable;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_6 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(global_clock_enable),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_6 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_hnj_5 auto_generated(
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clken(clken),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.result_i_tmp_8(result_i_tmp_8),
	.result_i_tmp_7(result_i_tmp_7),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.result_i_tmp_19(result_i_tmp_19),
	.result_i_tmp_18(result_i_tmp_18),
	.result_i_tmp_17(result_i_tmp_17),
	.result_i_tmp_16(result_i_tmp_16),
	.clock(clock));

endmodule

module fftsign_add_sub_hnj_5 (
	pipeline_dffe_15,
	pipeline_dffe_19,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_14,
	pipeline_dffe_13,
	clken,
	result_i_tmp_15,
	result_i_tmp_14,
	result_i_tmp_13,
	result_i_tmp_12,
	result_i_tmp_11,
	result_i_tmp_10,
	result_i_tmp_9,
	result_i_tmp_8,
	result_i_tmp_7,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	result_i_tmp_19,
	result_i_tmp_18,
	result_i_tmp_17,
	result_i_tmp_16,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_15;
output 	pipeline_dffe_19;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	clken;
input 	result_i_tmp_15;
input 	result_i_tmp_14;
input 	result_i_tmp_13;
input 	result_i_tmp_12;
input 	result_i_tmp_11;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
input 	result_i_tmp_8;
input 	result_i_tmp_7;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	result_i_tmp_19;
input 	result_i_tmp_18;
input 	result_i_tmp_17;
input 	result_i_tmp_16;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 (
	.dataa(result_i_tmp_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 (
	.dataa(result_i_tmp_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 (
	.dataa(result_i_tmp_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~15_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 (
	.dataa(result_i_tmp_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~17_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 (
	.dataa(result_i_tmp_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~19_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 (
	.dataa(result_i_tmp_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~21_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 (
	.dataa(result_i_tmp_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~23_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 (
	.dataa(result_i_tmp_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~25_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 (
	.dataa(result_i_tmp_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~27_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 (
	.dataa(result_i_tmp_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~29_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(result_i_tmp_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~31_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(result_i_tmp_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 (
	.dataa(result_i_tmp_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~35 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 (
	.dataa(result_i_tmp_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~37 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 (
	.dataa(result_i_tmp_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~39 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 (
	.dataa(result_i_tmp_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~41 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 (
	.dataa(result_i_tmp_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~43 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 (
	.dataa(result_i_tmp_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[16]~45 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 (
	.dataa(result_i_tmp_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[17]~47 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 (
	.dataa(result_i_tmp_19),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[18]~49 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_da0:gen_std:cm3|gen_ma:gen_ma_full:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[19]~50 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_tdl_4 (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_tdl_5 (
	data_in,
	global_clock_enable,
	tdl_arr_5_1,
	tdl_arr_9_1,
	tdl_arr_6_1,
	tdl_arr_7_1,
	tdl_arr_8_1,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	tdl_arr_4_1,
	tdl_arr_3_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_in;
input 	global_clock_enable;
output 	tdl_arr_5_1;
output 	tdl_arr_9_1;
output 	tdl_arr_6_1;
output 	tdl_arr_7_1;
output 	tdl_arr_8_1;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
output 	tdl_arr_4_1;
output 	tdl_arr_3_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][9]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][8]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][3]~q ;


dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][9] (
	.clk(clk),
	.d(\tdl_arr[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9_1),
	.prn(vcc));
defparam \tdl_arr[1][9] .is_wysiwyg = "true";
defparam \tdl_arr[1][9] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][8] (
	.clk(clk),
	.d(\tdl_arr[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_8_1),
	.prn(vcc));
defparam \tdl_arr[1][8] .is_wysiwyg = "true";
defparam \tdl_arr[1][8] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][9] (
	.clk(clk),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][9]~q ),
	.prn(vcc));
defparam \tdl_arr[0][9] .is_wysiwyg = "true";
defparam \tdl_arr[0][9] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][8] (
	.clk(clk),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][8]~q ),
	.prn(vcc));
defparam \tdl_arr[0][8] .is_wysiwyg = "true";
defparam \tdl_arr[0][8] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

endmodule

module fftsign_asj_fft_pround_6 (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2008,
	butterfly_st2007,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st20011,
	butterfly_st20010,
	butterfly_st2009,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st20011;
input 	butterfly_st20010;
input 	butterfly_st2009;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_7 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2007(butterfly_st2007),
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.butterfly_st20011(butterfly_st20011),
	.butterfly_st20010(butterfly_st20010),
	.butterfly_st2009(butterfly_st2009),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_7 (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2008,
	butterfly_st2007,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st20011,
	butterfly_st20010,
	butterfly_st2009,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st20011;
input 	butterfly_st20010;
input 	butterfly_st2009;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj auto_generated(
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2007(butterfly_st2007),
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.butterfly_st20011(butterfly_st20011),
	.butterfly_st20010(butterfly_st20010),
	.butterfly_st2009(butterfly_st2009),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2008,
	butterfly_st2007,
	butterfly_st2006,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	butterfly_st20011,
	butterfly_st20010,
	butterfly_st2009,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2008;
input 	butterfly_st2007;
input 	butterfly_st2006;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	butterfly_st20011;
input 	butterfly_st20010;
input 	butterfly_st2009;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st20011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2000),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2001),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2002),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2003),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2004),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2005),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2006),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2007),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2008),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2009),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st20010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st20011),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_7 (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	butterfly_st20111,
	butterfly_st20110,
	butterfly_st2019,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	butterfly_st20111;
input 	butterfly_st20110;
input 	butterfly_st2019;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_8 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.butterfly_st20111(butterfly_st20111),
	.butterfly_st20110(butterfly_st20110),
	.butterfly_st2019(butterfly_st2019),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_8 (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	butterfly_st20111,
	butterfly_st20110,
	butterfly_st2019,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	butterfly_st20111;
input 	butterfly_st20110;
input 	butterfly_st2019;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_1 auto_generated(
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.butterfly_st20111(butterfly_st20111),
	.butterfly_st20110(butterfly_st20110),
	.butterfly_st2019(butterfly_st2019),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_1 (
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	butterfly_st2018,
	butterfly_st2017,
	butterfly_st2016,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	butterfly_st20111,
	butterfly_st20110,
	butterfly_st2019,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
input 	butterfly_st2018;
input 	butterfly_st2017;
input 	butterfly_st2016;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	butterfly_st20111;
input 	butterfly_st20110;
input 	butterfly_st2019;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st20111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2012),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2013),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2014),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2015),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2016),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2017),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2018),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2019),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st20110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st20111),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_8 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st21011,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st21010,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st21011;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st21010;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_9 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.butterfly_st21011(butterfly_st21011),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st21010(butterfly_st21010),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st21011,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st21010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st21011;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st21010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_2 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.butterfly_st21011(butterfly_st21011),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st21010(butterfly_st21010),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_2 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2102,
	butterfly_st2101,
	butterfly_st2100,
	butterfly_st21011,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st21010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2102;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	butterfly_st21011;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st21010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st21011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2100),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2101),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2102),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2103),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2104),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2105),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2106),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2107),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2108),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2109),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st21010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st21011),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st21111,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st21110,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st21111;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st21110;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_10 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.butterfly_st21111(butterfly_st21111),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st21110(butterfly_st21110),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st21111,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st21110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st21111;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st21110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_3 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.butterfly_st21111(butterfly_st21111),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st21110(butterfly_st21110),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_3 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2112,
	butterfly_st2111,
	butterfly_st2110,
	butterfly_st21111,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st21110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2112;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	butterfly_st21111;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st21110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st21111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2112),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2113),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2114),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2115),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2116),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2117),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2118),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2119),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st21110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st21111),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st22011,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st22010,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st22011;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st22010;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_11 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.butterfly_st22011(butterfly_st22011),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st22010(butterfly_st22010),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st22011,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st22010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st22011;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st22010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_4 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.butterfly_st22011(butterfly_st22011),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st22010(butterfly_st22010),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_4 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2202,
	butterfly_st2201,
	butterfly_st2200,
	butterfly_st22011,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st22010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2202;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	butterfly_st22011;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st22010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st22011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2200),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2201),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2202),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2203),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2204),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2205),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2206),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2207),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2208),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2209),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st22010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st22011),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st22111,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st22110,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st22111;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st22110;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_12 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.butterfly_st22111(butterfly_st22111),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st22110(butterfly_st22110),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_12 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st22111,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st22110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st22111;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st22110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_5 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.butterfly_st22111(butterfly_st22111),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st22110(butterfly_st22110),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_5 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2212,
	butterfly_st2211,
	butterfly_st2210,
	butterfly_st22111,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st22110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2212;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	butterfly_st22111;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st22110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st22111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2210),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2211),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2212),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2213),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2214),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2215),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2216),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2217),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2218),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2219),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st22110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st22111),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_12 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st23011,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st23010,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st23011;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st23010;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_13 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.butterfly_st23011(butterfly_st23011),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st23010(butterfly_st23010),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_13 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st23011,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st23010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st23011;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st23010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_6 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.butterfly_st23011(butterfly_st23011),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st23010(butterfly_st23010),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_6 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2302,
	butterfly_st2301,
	butterfly_st2300,
	butterfly_st23011,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st23010,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2302;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	butterfly_st23011;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st23010;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st23011),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2300),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2301),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2302),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2303),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2304),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2305),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2306),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2307),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2308),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2309),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st23010),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st23011),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_13 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st23111,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st23110,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st23111;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st23110;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_14 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.butterfly_st23111(butterfly_st23111),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st23110(butterfly_st23110),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_14 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st23111,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st23110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st23111;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st23110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_7 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.butterfly_st23111(butterfly_st23111),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st23110(butterfly_st23110),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_7 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	butterfly_st2312,
	butterfly_st2311,
	butterfly_st2310,
	butterfly_st23111,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st23110,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	butterfly_st2312;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	butterfly_st23111;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st23110;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(butterfly_st23111),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(butterfly_st2310),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(butterfly_st2311),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(butterfly_st2312),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(butterfly_st2313),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(butterfly_st2314),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(butterfly_st2315),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(butterfly_st2316),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(butterfly_st2317),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(butterfly_st2318),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(butterfly_st2319),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(butterfly_st23110),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(butterfly_st23111),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_in_write_sgl (
	rdy_for_next_block1,
	disable_wr1,
	data_rdy_int1,
	wren_3,
	wren_0,
	wren_1,
	wren_2,
	blk_done_int,
	core_real_in_2,
	core_imag_in_2,
	core_real_in_1,
	core_imag_in_1,
	core_real_in_0,
	core_imag_in_0,
	core_real_in_9,
	core_imag_in_9,
	core_real_in_8,
	core_imag_in_8,
	core_real_in_7,
	core_imag_in_7,
	core_real_in_6,
	core_imag_in_6,
	core_real_in_5,
	core_imag_in_5,
	core_real_in_4,
	core_imag_in_4,
	core_real_in_3,
	core_imag_in_3,
	send_sop_s,
	global_clock_enable,
	data_in_r_2,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	wr_address_i_int_4,
	wr_address_i_int_5,
	wr_address_i_int_6,
	wr_address_i_int_7,
	data_in_i_2,
	data_in_r_1,
	data_in_i_1,
	data_in_r_0,
	data_in_i_0,
	data_in_r_9,
	data_in_i_9,
	data_in_r_8,
	data_in_i_8,
	data_in_r_7,
	data_in_i_7,
	data_in_r_6,
	data_in_i_6,
	data_in_r_5,
	data_in_i_5,
	data_in_r_4,
	data_in_i_4,
	data_in_r_3,
	data_in_i_3,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rdy_for_next_block1;
output 	disable_wr1;
output 	data_rdy_int1;
output 	wren_3;
output 	wren_0;
output 	wren_1;
output 	wren_2;
input 	blk_done_int;
input 	core_real_in_2;
input 	core_imag_in_2;
input 	core_real_in_1;
input 	core_imag_in_1;
input 	core_real_in_0;
input 	core_imag_in_0;
input 	core_real_in_9;
input 	core_imag_in_9;
input 	core_real_in_8;
input 	core_imag_in_8;
input 	core_real_in_7;
input 	core_imag_in_7;
input 	core_real_in_6;
input 	core_imag_in_6;
input 	core_real_in_5;
input 	core_imag_in_5;
input 	core_real_in_4;
input 	core_imag_in_4;
input 	core_real_in_3;
input 	core_imag_in_3;
input 	send_sop_s;
input 	global_clock_enable;
output 	data_in_r_2;
output 	wr_address_i_int_0;
output 	wr_address_i_int_1;
output 	wr_address_i_int_2;
output 	wr_address_i_int_3;
output 	wr_address_i_int_4;
output 	wr_address_i_int_5;
output 	wr_address_i_int_6;
output 	wr_address_i_int_7;
output 	data_in_i_2;
output 	data_in_r_1;
output 	data_in_i_1;
output 	data_in_r_0;
output 	data_in_i_0;
output 	data_in_r_9;
output 	data_in_i_9;
output 	data_in_r_8;
output 	data_in_i_8;
output 	data_in_r_7;
output 	data_in_i_7;
output 	data_in_r_6;
output 	data_in_i_6;
output 	data_in_r_5;
output 	data_in_i_5;
output 	data_in_r_4;
output 	data_in_i_4;
output 	data_in_r_3;
output 	data_in_i_3;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_quad:gen_se_writer:gen_burst_rdy:delay_swd|tdl_arr[0]~q ;
wire \count[0]~10_combout ;
wire \counter_i~0_combout ;
wire \burst_count_en~0_combout ;
wire \burst_count_en~q ;
wire \count[0]~16_combout ;
wire \count[0]~q ;
wire \count[0]~11 ;
wire \count[1]~12_combout ;
wire \count[1]~q ;
wire \count[1]~13 ;
wire \count[2]~14_combout ;
wire \count[2]~q ;
wire \count[2]~15 ;
wire \count[3]~17_combout ;
wire \count[3]~q ;
wire \count[3]~18 ;
wire \count[4]~19_combout ;
wire \count[4]~q ;
wire \count[4]~20 ;
wire \count[5]~21_combout ;
wire \count[5]~q ;
wire \count[5]~22 ;
wire \count[6]~23_combout ;
wire \count[6]~q ;
wire \count[6]~24 ;
wire \count[7]~25_combout ;
wire \count[7]~q ;
wire \count[7]~26 ;
wire \count[8]~27_combout ;
wire \count[8]~q ;
wire \Equal0~0_combout ;
wire \count[8]~28 ;
wire \count[9]~29_combout ;
wire \count[9]~q ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal1~0_combout ;
wire \data_rdy_int~0_combout ;
wire \Add1~0_combout ;
wire \sw[0]~q ;
wire \Add1~1_combout ;
wire \sw[1]~q ;
wire \Mux1~0_combout ;
wire \Mux3~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \data_in_r~0_combout ;
wire \wr_addr[0]~q ;
wire \wr_address_i_int~0_combout ;
wire \wr_addr[1]~q ;
wire \wr_address_i_int~1_combout ;
wire \wr_addr[2]~q ;
wire \wr_address_i_int~2_combout ;
wire \wr_addr[3]~q ;
wire \wr_address_i_int~3_combout ;
wire \wr_addr[4]~q ;
wire \wr_address_i_int~4_combout ;
wire \wr_addr[5]~q ;
wire \wr_address_i_int~5_combout ;
wire \wr_addr[6]~q ;
wire \wr_address_i_int~6_combout ;
wire \wr_addr[7]~q ;
wire \wr_address_i_int~7_combout ;
wire \data_in_i~0_combout ;
wire \data_in_r~1_combout ;
wire \data_in_i~1_combout ;
wire \data_in_r~2_combout ;
wire \data_in_i~2_combout ;
wire \data_in_r~3_combout ;
wire \data_in_i~3_combout ;
wire \data_in_r~4_combout ;
wire \data_in_i~4_combout ;
wire \data_in_r~5_combout ;
wire \data_in_i~5_combout ;
wire \data_in_r~6_combout ;
wire \data_in_i~6_combout ;
wire \data_in_r~7_combout ;
wire \data_in_i~7_combout ;
wire \data_in_r~8_combout ;
wire \data_in_i~8_combout ;
wire \data_in_r~9_combout ;
wire \data_in_i~9_combout ;


fftsign_asj_fft_tdl_bit_rst_3 \gen_quad:gen_se_writer:gen_burst_rdy:delay_swd (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0(\gen_quad:gen_se_writer:gen_burst_rdy:delay_swd|tdl_arr[0]~q ),
	.clk(clk),
	.reset_n(reset_n));

dffeas rdy_for_next_block(
	.clk(clk),
	.d(\Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdy_for_next_block1),
	.prn(vcc));
defparam rdy_for_next_block.is_wysiwyg = "true";
defparam rdy_for_next_block.power_up = "low";

dffeas disable_wr(
	.clk(clk),
	.d(\Equal1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(disable_wr1),
	.prn(vcc));
defparam disable_wr.is_wysiwyg = "true";
defparam disable_wr.power_up = "low";

dffeas data_rdy_int(
	.clk(clk),
	.d(\data_rdy_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_rdy_int1),
	.prn(vcc));
defparam data_rdy_int.is_wysiwyg = "true";
defparam data_rdy_int.power_up = "low";

dffeas \wren[3] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_3),
	.prn(vcc));
defparam \wren[3] .is_wysiwyg = "true";
defparam \wren[3] .power_up = "low";

dffeas \wren[0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_0),
	.prn(vcc));
defparam \wren[0] .is_wysiwyg = "true";
defparam \wren[0] .power_up = "low";

dffeas \wren[1] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_1),
	.prn(vcc));
defparam \wren[1] .is_wysiwyg = "true";
defparam \wren[1] .power_up = "low";

dffeas \wren[2] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wren_2),
	.prn(vcc));
defparam \wren[2] .is_wysiwyg = "true";
defparam \wren[2] .power_up = "low";

dffeas \data_in_r[2] (
	.clk(clk),
	.d(\data_in_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_2),
	.prn(vcc));
defparam \data_in_r[2] .is_wysiwyg = "true";
defparam \data_in_r[2] .power_up = "low";

dffeas \wr_address_i_int[0] (
	.clk(clk),
	.d(\wr_address_i_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_0),
	.prn(vcc));
defparam \wr_address_i_int[0] .is_wysiwyg = "true";
defparam \wr_address_i_int[0] .power_up = "low";

dffeas \wr_address_i_int[1] (
	.clk(clk),
	.d(\wr_address_i_int~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_1),
	.prn(vcc));
defparam \wr_address_i_int[1] .is_wysiwyg = "true";
defparam \wr_address_i_int[1] .power_up = "low";

dffeas \wr_address_i_int[2] (
	.clk(clk),
	.d(\wr_address_i_int~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_2),
	.prn(vcc));
defparam \wr_address_i_int[2] .is_wysiwyg = "true";
defparam \wr_address_i_int[2] .power_up = "low";

dffeas \wr_address_i_int[3] (
	.clk(clk),
	.d(\wr_address_i_int~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_3),
	.prn(vcc));
defparam \wr_address_i_int[3] .is_wysiwyg = "true";
defparam \wr_address_i_int[3] .power_up = "low";

dffeas \wr_address_i_int[4] (
	.clk(clk),
	.d(\wr_address_i_int~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_4),
	.prn(vcc));
defparam \wr_address_i_int[4] .is_wysiwyg = "true";
defparam \wr_address_i_int[4] .power_up = "low";

dffeas \wr_address_i_int[5] (
	.clk(clk),
	.d(\wr_address_i_int~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_5),
	.prn(vcc));
defparam \wr_address_i_int[5] .is_wysiwyg = "true";
defparam \wr_address_i_int[5] .power_up = "low";

dffeas \wr_address_i_int[6] (
	.clk(clk),
	.d(\wr_address_i_int~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_6),
	.prn(vcc));
defparam \wr_address_i_int[6] .is_wysiwyg = "true";
defparam \wr_address_i_int[6] .power_up = "low";

dffeas \wr_address_i_int[7] (
	.clk(clk),
	.d(\wr_address_i_int~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wr_address_i_int_7),
	.prn(vcc));
defparam \wr_address_i_int[7] .is_wysiwyg = "true";
defparam \wr_address_i_int[7] .power_up = "low";

dffeas \data_in_i[2] (
	.clk(clk),
	.d(\data_in_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_2),
	.prn(vcc));
defparam \data_in_i[2] .is_wysiwyg = "true";
defparam \data_in_i[2] .power_up = "low";

dffeas \data_in_r[1] (
	.clk(clk),
	.d(\data_in_r~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_1),
	.prn(vcc));
defparam \data_in_r[1] .is_wysiwyg = "true";
defparam \data_in_r[1] .power_up = "low";

dffeas \data_in_i[1] (
	.clk(clk),
	.d(\data_in_i~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_1),
	.prn(vcc));
defparam \data_in_i[1] .is_wysiwyg = "true";
defparam \data_in_i[1] .power_up = "low";

dffeas \data_in_r[0] (
	.clk(clk),
	.d(\data_in_r~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_0),
	.prn(vcc));
defparam \data_in_r[0] .is_wysiwyg = "true";
defparam \data_in_r[0] .power_up = "low";

dffeas \data_in_i[0] (
	.clk(clk),
	.d(\data_in_i~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_0),
	.prn(vcc));
defparam \data_in_i[0] .is_wysiwyg = "true";
defparam \data_in_i[0] .power_up = "low";

dffeas \data_in_r[9] (
	.clk(clk),
	.d(\data_in_r~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_9),
	.prn(vcc));
defparam \data_in_r[9] .is_wysiwyg = "true";
defparam \data_in_r[9] .power_up = "low";

dffeas \data_in_i[9] (
	.clk(clk),
	.d(\data_in_i~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_9),
	.prn(vcc));
defparam \data_in_i[9] .is_wysiwyg = "true";
defparam \data_in_i[9] .power_up = "low";

dffeas \data_in_r[8] (
	.clk(clk),
	.d(\data_in_r~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_8),
	.prn(vcc));
defparam \data_in_r[8] .is_wysiwyg = "true";
defparam \data_in_r[8] .power_up = "low";

dffeas \data_in_i[8] (
	.clk(clk),
	.d(\data_in_i~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_8),
	.prn(vcc));
defparam \data_in_i[8] .is_wysiwyg = "true";
defparam \data_in_i[8] .power_up = "low";

dffeas \data_in_r[7] (
	.clk(clk),
	.d(\data_in_r~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_7),
	.prn(vcc));
defparam \data_in_r[7] .is_wysiwyg = "true";
defparam \data_in_r[7] .power_up = "low";

dffeas \data_in_i[7] (
	.clk(clk),
	.d(\data_in_i~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_7),
	.prn(vcc));
defparam \data_in_i[7] .is_wysiwyg = "true";
defparam \data_in_i[7] .power_up = "low";

dffeas \data_in_r[6] (
	.clk(clk),
	.d(\data_in_r~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_6),
	.prn(vcc));
defparam \data_in_r[6] .is_wysiwyg = "true";
defparam \data_in_r[6] .power_up = "low";

dffeas \data_in_i[6] (
	.clk(clk),
	.d(\data_in_i~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_6),
	.prn(vcc));
defparam \data_in_i[6] .is_wysiwyg = "true";
defparam \data_in_i[6] .power_up = "low";

dffeas \data_in_r[5] (
	.clk(clk),
	.d(\data_in_r~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_5),
	.prn(vcc));
defparam \data_in_r[5] .is_wysiwyg = "true";
defparam \data_in_r[5] .power_up = "low";

dffeas \data_in_i[5] (
	.clk(clk),
	.d(\data_in_i~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_5),
	.prn(vcc));
defparam \data_in_i[5] .is_wysiwyg = "true";
defparam \data_in_i[5] .power_up = "low";

dffeas \data_in_r[4] (
	.clk(clk),
	.d(\data_in_r~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_4),
	.prn(vcc));
defparam \data_in_r[4] .is_wysiwyg = "true";
defparam \data_in_r[4] .power_up = "low";

dffeas \data_in_i[4] (
	.clk(clk),
	.d(\data_in_i~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_4),
	.prn(vcc));
defparam \data_in_i[4] .is_wysiwyg = "true";
defparam \data_in_i[4] .power_up = "low";

dffeas \data_in_r[3] (
	.clk(clk),
	.d(\data_in_r~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_r_3),
	.prn(vcc));
defparam \data_in_r[3] .is_wysiwyg = "true";
defparam \data_in_r[3] .power_up = "low";

dffeas \data_in_i[3] (
	.clk(clk),
	.d(\data_in_i~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_in_i_3),
	.prn(vcc));
defparam \data_in_i[3] .is_wysiwyg = "true";
defparam \data_in_i[3] .power_up = "low";

cycloneive_lcell_comb \count[0]~10 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~10_combout ),
	.cout(\count[0]~11 ));
defparam \count[0]~10 .lut_mask = 16'h55AA;
defparam \count[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \counter_i~0 (
	.dataa(send_sop_s),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\counter_i~0_combout ),
	.cout());
defparam \counter_i~0 .lut_mask = 16'hAAFF;
defparam \counter_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burst_count_en~0 (
	.dataa(send_sop_s),
	.datab(\burst_count_en~q ),
	.datac(gnd),
	.datad(rdy_for_next_block1),
	.cin(gnd),
	.combout(\burst_count_en~0_combout ),
	.cout());
defparam \burst_count_en~0 .lut_mask = 16'hEEFF;
defparam \burst_count_en~0 .sum_lutc_input = "datac";

dffeas burst_count_en(
	.clk(clk),
	.d(\burst_count_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\burst_count_en~q ),
	.prn(vcc));
defparam burst_count_en.is_wysiwyg = "true";
defparam burst_count_en.power_up = "low";

cycloneive_lcell_comb \count[0]~16 (
	.dataa(global_clock_enable),
	.datab(\gen_quad:gen_se_writer:gen_burst_rdy:delay_swd|tdl_arr[0]~q ),
	.datac(\burst_count_en~q ),
	.datad(\counter_i~0_combout ),
	.cin(gnd),
	.combout(\count[0]~16_combout ),
	.cout());
defparam \count[0]~16 .lut_mask = 16'hFFFE;
defparam \count[0]~16 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \count[1]~12 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~11 ),
	.combout(\count[1]~12_combout ),
	.cout(\count[1]~13 ));
defparam \count[1]~12 .lut_mask = 16'h5A5F;
defparam \count[1]~12 .sum_lutc_input = "cin";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \count[2]~14 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~13 ),
	.combout(\count[2]~14_combout ),
	.cout(\count[2]~15 ));
defparam \count[2]~14 .lut_mask = 16'h5AAF;
defparam \count[2]~14 .sum_lutc_input = "cin";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count[3]~17 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~15 ),
	.combout(\count[3]~17_combout ),
	.cout(\count[3]~18 ));
defparam \count[3]~17 .lut_mask = 16'h5A5F;
defparam \count[3]~17 .sum_lutc_input = "cin";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count[4]~19 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~18 ),
	.combout(\count[4]~19_combout ),
	.cout(\count[4]~20 ));
defparam \count[4]~19 .lut_mask = 16'h5AAF;
defparam \count[4]~19 .sum_lutc_input = "cin";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count[5]~21 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~20 ),
	.combout(\count[5]~21_combout ),
	.cout(\count[5]~22 ));
defparam \count[5]~21 .lut_mask = 16'h5A5F;
defparam \count[5]~21 .sum_lutc_input = "cin";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count[6]~23 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~22 ),
	.combout(\count[6]~23_combout ),
	.cout(\count[6]~24 ));
defparam \count[6]~23 .lut_mask = 16'h5AAF;
defparam \count[6]~23 .sum_lutc_input = "cin";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count[7]~25 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~24 ),
	.combout(\count[7]~25_combout ),
	.cout(\count[7]~26 ));
defparam \count[7]~25 .lut_mask = 16'h5A5F;
defparam \count[7]~25 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \count[8]~27 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[7]~26 ),
	.combout(\count[8]~27_combout ),
	.cout(\count[8]~28 ));
defparam \count[8]~27 .lut_mask = 16'h5AAF;
defparam \count[8]~27 .sum_lutc_input = "cin";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\count[0]~q ),
	.datab(\count[8]~q ),
	.datac(\count[1]~q ),
	.datad(\count[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[9]~29 (
	.dataa(\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[8]~28 ),
	.combout(\count[9]~29_combout ),
	.cout());
defparam \count[9]~29 .lut_mask = 16'h5A5A;
defparam \count[9]~29 .sum_lutc_input = "cin";

dffeas \count[9] (
	.clk(clk),
	.d(\count[9]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(\count[0]~16_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\count[4]~q ),
	.datab(\count[5]~q ),
	.datac(\count[6]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFFFE;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\count[2]~q ),
	.datab(\Equal0~0_combout ),
	.datac(\count[9]~q ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFFFE;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\Equal0~0_combout ),
	.datab(\count[9]~q ),
	.datac(\Equal0~1_combout ),
	.datad(\count[2]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_rdy_int~0 (
	.dataa(rdy_for_next_block1),
	.datab(data_rdy_int1),
	.datac(gnd),
	.datad(blk_done_int),
	.cin(gnd),
	.combout(\data_rdy_int~0_combout ),
	.cout());
defparam \data_rdy_int~0 .lut_mask = 16'hEEFF;
defparam \data_rdy_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\count[0]~q ),
	.datad(\count[8]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas \sw[0] (
	.clk(clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw[0]~q ),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\count[0]~q ),
	.datab(\count[8]~q ),
	.datac(\count[1]~q ),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

dffeas \sw[1] (
	.clk(clk),
	.d(\Add1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sw[1]~q ),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\sw[0]~q ),
	.datab(\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEEEE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\sw[0]~q ),
	.datab(\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'h7777;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(\sw[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sw[1]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hAAFF;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(\sw[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sw[0]~q ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hAAFF;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~0 (
	.dataa(reset_n),
	.datab(core_real_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~0_combout ),
	.cout());
defparam \data_in_r~0 .lut_mask = 16'hEEEE;
defparam \data_in_r~0 .sum_lutc_input = "datac";

dffeas \wr_addr[0] (
	.clk(clk),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[0]~q ),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~0 (
	.dataa(reset_n),
	.datab(\wr_addr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~0_combout ),
	.cout());
defparam \wr_address_i_int~0 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~0 .sum_lutc_input = "datac";

dffeas \wr_addr[1] (
	.clk(clk),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[1]~q ),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~1 (
	.dataa(reset_n),
	.datab(\wr_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~1_combout ),
	.cout());
defparam \wr_address_i_int~1 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~1 .sum_lutc_input = "datac";

dffeas \wr_addr[2] (
	.clk(clk),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[2]~q ),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~2 (
	.dataa(reset_n),
	.datab(\wr_addr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~2_combout ),
	.cout());
defparam \wr_address_i_int~2 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~2 .sum_lutc_input = "datac";

dffeas \wr_addr[3] (
	.clk(clk),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[3]~q ),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~3 (
	.dataa(reset_n),
	.datab(\wr_addr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~3_combout ),
	.cout());
defparam \wr_address_i_int~3 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~3 .sum_lutc_input = "datac";

dffeas \wr_addr[4] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[4]~q ),
	.prn(vcc));
defparam \wr_addr[4] .is_wysiwyg = "true";
defparam \wr_addr[4] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~4 (
	.dataa(reset_n),
	.datab(\wr_addr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~4_combout ),
	.cout());
defparam \wr_address_i_int~4 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~4 .sum_lutc_input = "datac";

dffeas \wr_addr[5] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[5]~q ),
	.prn(vcc));
defparam \wr_addr[5] .is_wysiwyg = "true";
defparam \wr_addr[5] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~5 (
	.dataa(reset_n),
	.datab(\wr_addr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~5_combout ),
	.cout());
defparam \wr_address_i_int~5 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~5 .sum_lutc_input = "datac";

dffeas \wr_addr[6] (
	.clk(clk),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[6]~q ),
	.prn(vcc));
defparam \wr_addr[6] .is_wysiwyg = "true";
defparam \wr_addr[6] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~6 (
	.dataa(reset_n),
	.datab(\wr_addr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~6_combout ),
	.cout());
defparam \wr_address_i_int~6 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~6 .sum_lutc_input = "datac";

dffeas \wr_addr[7] (
	.clk(clk),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\wr_addr[7]~q ),
	.prn(vcc));
defparam \wr_addr[7] .is_wysiwyg = "true";
defparam \wr_addr[7] .power_up = "low";

cycloneive_lcell_comb \wr_address_i_int~7 (
	.dataa(reset_n),
	.datab(\wr_addr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_address_i_int~7_combout ),
	.cout());
defparam \wr_address_i_int~7 .lut_mask = 16'hEEEE;
defparam \wr_address_i_int~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~0 (
	.dataa(reset_n),
	.datab(core_imag_in_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~0_combout ),
	.cout());
defparam \data_in_i~0 .lut_mask = 16'hEEEE;
defparam \data_in_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~1 (
	.dataa(reset_n),
	.datab(core_real_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~1_combout ),
	.cout());
defparam \data_in_r~1 .lut_mask = 16'hEEEE;
defparam \data_in_r~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~1 (
	.dataa(reset_n),
	.datab(core_imag_in_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~1_combout ),
	.cout());
defparam \data_in_i~1 .lut_mask = 16'hEEEE;
defparam \data_in_i~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~2 (
	.dataa(reset_n),
	.datab(core_real_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~2_combout ),
	.cout());
defparam \data_in_r~2 .lut_mask = 16'hEEEE;
defparam \data_in_r~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~2 (
	.dataa(reset_n),
	.datab(core_imag_in_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~2_combout ),
	.cout());
defparam \data_in_i~2 .lut_mask = 16'hEEEE;
defparam \data_in_i~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~3 (
	.dataa(reset_n),
	.datab(core_real_in_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~3_combout ),
	.cout());
defparam \data_in_r~3 .lut_mask = 16'hEEEE;
defparam \data_in_r~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~3 (
	.dataa(reset_n),
	.datab(core_imag_in_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~3_combout ),
	.cout());
defparam \data_in_i~3 .lut_mask = 16'hEEEE;
defparam \data_in_i~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~4 (
	.dataa(reset_n),
	.datab(core_real_in_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~4_combout ),
	.cout());
defparam \data_in_r~4 .lut_mask = 16'hEEEE;
defparam \data_in_r~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~4 (
	.dataa(reset_n),
	.datab(core_imag_in_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~4_combout ),
	.cout());
defparam \data_in_i~4 .lut_mask = 16'hEEEE;
defparam \data_in_i~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~5 (
	.dataa(reset_n),
	.datab(core_real_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~5_combout ),
	.cout());
defparam \data_in_r~5 .lut_mask = 16'hEEEE;
defparam \data_in_r~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~5 (
	.dataa(reset_n),
	.datab(core_imag_in_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~5_combout ),
	.cout());
defparam \data_in_i~5 .lut_mask = 16'hEEEE;
defparam \data_in_i~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~6 (
	.dataa(reset_n),
	.datab(core_real_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~6_combout ),
	.cout());
defparam \data_in_r~6 .lut_mask = 16'hEEEE;
defparam \data_in_r~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~6 (
	.dataa(reset_n),
	.datab(core_imag_in_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~6_combout ),
	.cout());
defparam \data_in_i~6 .lut_mask = 16'hEEEE;
defparam \data_in_i~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~7 (
	.dataa(reset_n),
	.datab(core_real_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~7_combout ),
	.cout());
defparam \data_in_r~7 .lut_mask = 16'hEEEE;
defparam \data_in_r~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~7 (
	.dataa(reset_n),
	.datab(core_imag_in_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~7_combout ),
	.cout());
defparam \data_in_i~7 .lut_mask = 16'hEEEE;
defparam \data_in_i~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~8 (
	.dataa(reset_n),
	.datab(core_real_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~8_combout ),
	.cout());
defparam \data_in_r~8 .lut_mask = 16'hEEEE;
defparam \data_in_r~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~8 (
	.dataa(reset_n),
	.datab(core_imag_in_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~8_combout ),
	.cout());
defparam \data_in_i~8 .lut_mask = 16'hEEEE;
defparam \data_in_i~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_r~9 (
	.dataa(reset_n),
	.datab(core_real_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_r~9_combout ),
	.cout());
defparam \data_in_r~9 .lut_mask = 16'hEEEE;
defparam \data_in_r~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_i~9 (
	.dataa(reset_n),
	.datab(core_imag_in_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_in_i~9_combout ),
	.cout());
defparam \data_in_i~9 .lut_mask = 16'hEEEE;
defparam \data_in_i~9 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_rst_3 (
	global_clock_enable,
	tdl_arr_0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module fftsign_asj_fft_lpp_serial (
	ram_in_reg_2_3,
	ram_in_reg_2_7,
	ram_in_reg_2_1,
	ram_in_reg_2_5,
	ram_in_reg_1_3,
	ram_in_reg_1_7,
	ram_in_reg_1_1,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	ram_in_reg_0_1,
	ram_in_reg_0_5,
	data_3_imag_i,
	data_1_imag_i,
	ram_in_reg_9_3,
	ram_in_reg_9_7,
	ram_in_reg_9_1,
	ram_in_reg_9_5,
	ram_in_reg_8_3,
	ram_in_reg_8_7,
	ram_in_reg_8_1,
	ram_in_reg_8_5,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	data_3_real_i,
	data_1_real_i,
	global_clock_enable,
	data_imag_o_0,
	data_real_o_0,
	data_imag_o_1,
	data_real_o_1,
	data_imag_o_2,
	data_real_o_2,
	data_imag_o_3,
	data_real_o_3,
	data_imag_o_4,
	data_real_o_4,
	data_imag_o_5,
	data_real_o_5,
	data_imag_o_6,
	data_real_o_6,
	data_imag_o_7,
	data_real_o_7,
	data_imag_o_8,
	data_real_o_8,
	data_imag_o_9,
	data_real_o_9,
	wait_count_0,
	tdl_arr_4,
	tdl_arr_41,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	ram_in_reg_2_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_1;
input 	ram_in_reg_2_5;
input 	ram_in_reg_1_3;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_5;
input 	[9:0] data_3_imag_i;
input 	[9:0] data_1_imag_i;
input 	ram_in_reg_9_3;
input 	ram_in_reg_9_7;
input 	ram_in_reg_9_1;
input 	ram_in_reg_9_5;
input 	ram_in_reg_8_3;
input 	ram_in_reg_8_7;
input 	ram_in_reg_8_1;
input 	ram_in_reg_8_5;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	[9:0] data_3_real_i;
input 	[9:0] data_1_real_i;
input 	global_clock_enable;
output 	data_imag_o_0;
output 	data_real_o_0;
output 	data_imag_o_1;
output 	data_real_o_1;
output 	data_imag_o_2;
output 	data_real_o_2;
output 	data_imag_o_3;
output 	data_real_o_3;
output 	data_imag_o_4;
output 	data_real_o_4;
output 	data_imag_o_5;
output 	data_real_o_5;
output 	data_imag_o_6;
output 	data_real_o_6;
output 	data_imag_o_7;
output 	data_real_o_7;
output 	data_imag_o_8;
output 	data_real_o_8;
output 	data_imag_o_9;
output 	data_real_o_9;
input 	wait_count_0;
input 	tdl_arr_4;
output 	tdl_arr_41;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \output_i[2]~q ;
wire \output_i[1]~q ;
wire \output_i[0]~q ;
wire \output_i[11]~q ;
wire \output_r[2]~q ;
wire \output_r[1]~q ;
wire \output_r[0]~q ;
wire \output_r[11]~q ;
wire \output_i[3]~q ;
wire \output_r[3]~q ;
wire \output_i[4]~q ;
wire \output_r[4]~q ;
wire \output_i[5]~q ;
wire \output_r[5]~q ;
wire \output_i[6]~q ;
wire \output_r[6]~q ;
wire \output_i[7]~q ;
wire \output_r[7]~q ;
wire \output_i[8]~q ;
wire \output_r[8]~q ;
wire \output_i[9]~q ;
wire \output_r[9]~q ;
wire \output_i[10]~q ;
wire \output_r[10]~q ;
wire \result_ib[2]~q ;
wire \result_ia[2]~q ;
wire \result_ib[1]~q ;
wire \result_ia[1]~q ;
wire \result_ib[0]~q ;
wire \result_ia[0]~q ;
wire \output_i[0]~13_cout ;
wire \output_i[0]~15 ;
wire \output_i[0]~14_combout ;
wire \output_i[1]~17 ;
wire \output_i[1]~16_combout ;
wire \output_i[2]~19 ;
wire \output_i[2]~18_combout ;
wire \result_ib[10]~q ;
wire \result_ia[10]~q ;
wire \result_ib[9]~q ;
wire \result_ia[9]~q ;
wire \result_ib[8]~q ;
wire \result_ia[8]~q ;
wire \result_ib[7]~q ;
wire \result_ia[7]~q ;
wire \result_ib[6]~q ;
wire \result_ia[6]~q ;
wire \result_ib[5]~q ;
wire \result_ia[5]~q ;
wire \result_ib[4]~q ;
wire \result_ia[4]~q ;
wire \result_ib[3]~q ;
wire \result_ia[3]~q ;
wire \output_i[3]~21 ;
wire \output_i[3]~20_combout ;
wire \output_i[4]~23 ;
wire \output_i[4]~22_combout ;
wire \output_i[5]~25 ;
wire \output_i[5]~24_combout ;
wire \output_i[6]~27 ;
wire \output_i[6]~26_combout ;
wire \output_i[7]~29 ;
wire \output_i[7]~28_combout ;
wire \output_i[8]~31 ;
wire \output_i[8]~30_combout ;
wire \output_i[9]~33 ;
wire \output_i[9]~32_combout ;
wire \output_i[10]~35 ;
wire \output_i[10]~34_combout ;
wire \output_i[11]~36_combout ;
wire \result_rb[2]~q ;
wire \result_ra[2]~q ;
wire \result_rb[1]~q ;
wire \result_ra[1]~q ;
wire \result_rb[0]~q ;
wire \result_ra[0]~q ;
wire \output_r[0]~13_cout ;
wire \output_r[0]~15 ;
wire \output_r[0]~14_combout ;
wire \output_r[1]~17 ;
wire \output_r[1]~16_combout ;
wire \output_r[2]~19 ;
wire \output_r[2]~18_combout ;
wire \result_rb[10]~q ;
wire \result_ra[10]~q ;
wire \result_rb[9]~q ;
wire \result_ra[9]~q ;
wire \result_rb[8]~q ;
wire \result_ra[8]~q ;
wire \result_rb[7]~q ;
wire \result_ra[7]~q ;
wire \result_rb[6]~q ;
wire \result_ra[6]~q ;
wire \result_rb[5]~q ;
wire \result_ra[5]~q ;
wire \result_rb[4]~q ;
wire \result_ra[4]~q ;
wire \result_rb[3]~q ;
wire \result_ra[3]~q ;
wire \output_r[3]~21 ;
wire \output_r[3]~20_combout ;
wire \output_r[4]~23 ;
wire \output_r[4]~22_combout ;
wire \output_r[5]~25 ;
wire \output_r[5]~24_combout ;
wire \output_r[6]~27 ;
wire \output_r[6]~26_combout ;
wire \output_r[7]~29 ;
wire \output_r[7]~28_combout ;
wire \output_r[8]~31 ;
wire \output_r[8]~30_combout ;
wire \output_r[9]~33 ;
wire \output_r[9]~32_combout ;
wire \output_r[10]~35 ;
wire \output_r[10]~34_combout ;
wire \output_r[11]~36_combout ;
wire \result_ib[0]~12_cout ;
wire \result_ib[0]~14 ;
wire \result_ib[0]~13_combout ;
wire \result_ib[1]~16 ;
wire \result_ib[1]~15_combout ;
wire \result_ib[2]~18 ;
wire \result_ib[2]~17_combout ;
wire \result_ia[0]~12_cout ;
wire \result_ia[0]~14 ;
wire \result_ia[0]~13_combout ;
wire \result_ia[1]~16 ;
wire \result_ia[1]~15_combout ;
wire \result_ia[2]~18 ;
wire \result_ia[2]~17_combout ;
wire \result_ib[3]~20 ;
wire \result_ib[3]~19_combout ;
wire \result_ib[4]~22 ;
wire \result_ib[4]~21_combout ;
wire \result_ib[5]~24 ;
wire \result_ib[5]~23_combout ;
wire \result_ib[6]~26 ;
wire \result_ib[6]~25_combout ;
wire \result_ib[7]~28 ;
wire \result_ib[7]~27_combout ;
wire \result_ib[8]~30 ;
wire \result_ib[8]~29_combout ;
wire \result_ib[9]~32 ;
wire \result_ib[9]~31_combout ;
wire \result_ib[10]~33_combout ;
wire \result_ia[3]~20 ;
wire \result_ia[3]~19_combout ;
wire \result_ia[4]~22 ;
wire \result_ia[4]~21_combout ;
wire \result_ia[5]~24 ;
wire \result_ia[5]~23_combout ;
wire \result_ia[6]~26 ;
wire \result_ia[6]~25_combout ;
wire \result_ia[7]~28 ;
wire \result_ia[7]~27_combout ;
wire \result_ia[8]~30 ;
wire \result_ia[8]~29_combout ;
wire \result_ia[9]~32 ;
wire \result_ia[9]~31_combout ;
wire \result_ia[10]~33_combout ;
wire \result_rb[0]~12_cout ;
wire \result_rb[0]~14 ;
wire \result_rb[0]~13_combout ;
wire \result_rb[1]~16 ;
wire \result_rb[1]~15_combout ;
wire \result_rb[2]~18 ;
wire \result_rb[2]~17_combout ;
wire \result_ra[0]~12_cout ;
wire \result_ra[0]~14 ;
wire \result_ra[0]~13_combout ;
wire \result_ra[1]~16 ;
wire \result_ra[1]~15_combout ;
wire \result_ra[2]~18 ;
wire \result_ra[2]~17_combout ;
wire \result_rb[3]~20 ;
wire \result_rb[3]~19_combout ;
wire \result_rb[4]~22 ;
wire \result_rb[4]~21_combout ;
wire \result_rb[5]~24 ;
wire \result_rb[5]~23_combout ;
wire \result_rb[6]~26 ;
wire \result_rb[6]~25_combout ;
wire \result_rb[7]~28 ;
wire \result_rb[7]~27_combout ;
wire \result_rb[8]~30 ;
wire \result_rb[8]~29_combout ;
wire \result_rb[9]~32 ;
wire \result_rb[9]~31_combout ;
wire \result_rb[10]~33_combout ;
wire \result_ra[3]~20 ;
wire \result_ra[3]~19_combout ;
wire \result_ra[4]~22 ;
wire \result_ra[4]~21_combout ;
wire \result_ra[5]~24 ;
wire \result_ra[5]~23_combout ;
wire \result_ra[6]~26 ;
wire \result_ra[6]~25_combout ;
wire \result_ra[7]~28 ;
wire \result_ra[7]~27_combout ;
wire \result_ra[8]~30 ;
wire \result_ra[8]~29_combout ;
wire \result_ra[9]~32 ;
wire \result_ra[9]~31_combout ;
wire \result_ra[10]~33_combout ;
wire \offset_counter[8]~q ;
wire \offset_counter[9]~q ;
wire \data_val_i~q ;
wire \offset_counter[7]~q ;
wire \offset_counter[6]~q ;
wire \offset_counter[5]~q ;
wire \offset_counter[4]~q ;
wire \offset_counter[3]~q ;
wire \offset_counter[2]~q ;
wire \offset_counter[1]~q ;
wire \offset_counter[0]~q ;
wire \offset_counter[0]~11 ;
wire \offset_counter[0]~10_combout ;
wire \offset_counter[1]~13 ;
wire \offset_counter[1]~12_combout ;
wire \offset_counter[2]~15 ;
wire \offset_counter[2]~14_combout ;
wire \offset_counter[3]~17 ;
wire \offset_counter[3]~16_combout ;
wire \offset_counter[4]~19 ;
wire \offset_counter[4]~18_combout ;
wire \offset_counter[5]~21 ;
wire \offset_counter[5]~20_combout ;
wire \offset_counter[6]~23 ;
wire \offset_counter[6]~22_combout ;
wire \offset_counter[7]~25 ;
wire \offset_counter[7]~24_combout ;
wire \offset_counter[8]~27 ;
wire \offset_counter[8]~26_combout ;
wire \offset_counter[9]~29_combout ;
wire \sgn_2i~q ;
wire \Add11~0_combout ;
wire \Add11~1_combout ;
wire \Add11~2_combout ;
wire \Add11~3_combout ;
wire \Add11~4_combout ;
wire \Add11~5_combout ;
wire \Add11~6_combout ;
wire \Add11~7_combout ;
wire \Add11~8_combout ;
wire \Add11~9_combout ;
wire \Add11~10_combout ;
wire \sgn_2r~q ;
wire \Add9~0_combout ;
wire \Add9~1_combout ;
wire \Add9~2_combout ;
wire \Add9~3_combout ;
wire \Add9~4_combout ;
wire \Add9~5_combout ;
wire \Add9~6_combout ;
wire \Add9~7_combout ;
wire \Add9~8_combout ;
wire \Add9~9_combout ;
wire \Add9~10_combout ;
wire \sign_vec[0]~q ;
wire \add_in_i_d[2]~q ;
wire \sign_vec[3]~q ;
wire \Add4~0_combout ;
wire \add_in_i_c[2]~q ;
wire \add_in_i_d[1]~q ;
wire \Add4~1_combout ;
wire \add_in_i_c[1]~q ;
wire \add_in_i_d[0]~q ;
wire \Add4~2_combout ;
wire \add_in_i_c[0]~q ;
wire \add_in_i_b[2]~q ;
wire \Add2~0_combout ;
wire \add_in_i_a[2]~q ;
wire \add_in_i_b[1]~q ;
wire \Add2~1_combout ;
wire \add_in_i_a[1]~q ;
wire \add_in_i_b[0]~q ;
wire \Add2~2_combout ;
wire \add_in_i_a[0]~q ;
wire \add_in_i_d[9]~q ;
wire \Add4~3_combout ;
wire \add_in_i_c[9]~q ;
wire \add_in_i_d[8]~q ;
wire \Add4~4_combout ;
wire \add_in_i_c[8]~q ;
wire \add_in_i_d[7]~q ;
wire \Add4~5_combout ;
wire \add_in_i_c[7]~q ;
wire \add_in_i_d[6]~q ;
wire \Add4~6_combout ;
wire \add_in_i_c[6]~q ;
wire \add_in_i_d[5]~q ;
wire \Add4~7_combout ;
wire \add_in_i_c[5]~q ;
wire \add_in_i_d[4]~q ;
wire \Add4~8_combout ;
wire \add_in_i_c[4]~q ;
wire \add_in_i_d[3]~q ;
wire \Add4~9_combout ;
wire \add_in_i_c[3]~q ;
wire \add_in_i_b[9]~q ;
wire \Add2~3_combout ;
wire \add_in_i_a[9]~q ;
wire \add_in_i_b[8]~q ;
wire \Add2~4_combout ;
wire \add_in_i_a[8]~q ;
wire \add_in_i_b[7]~q ;
wire \Add2~5_combout ;
wire \add_in_i_a[7]~q ;
wire \add_in_i_b[6]~q ;
wire \Add2~6_combout ;
wire \add_in_i_a[6]~q ;
wire \add_in_i_b[5]~q ;
wire \Add2~7_combout ;
wire \add_in_i_a[5]~q ;
wire \add_in_i_b[4]~q ;
wire \Add2~8_combout ;
wire \add_in_i_a[4]~q ;
wire \add_in_i_b[3]~q ;
wire \Add2~9_combout ;
wire \add_in_i_a[3]~q ;
wire \sign_vec[1]~q ;
wire \add_in_r_d[2]~q ;
wire \Add3~0_combout ;
wire \add_in_r_c[2]~q ;
wire \add_in_r_d[1]~q ;
wire \Add3~1_combout ;
wire \add_in_r_c[1]~q ;
wire \add_in_r_d[0]~q ;
wire \Add3~2_combout ;
wire \add_in_r_c[0]~q ;
wire \add_in_r_b[2]~q ;
wire \Add1~0_combout ;
wire \add_in_r_a[2]~q ;
wire \add_in_r_b[1]~q ;
wire \Add1~1_combout ;
wire \add_in_r_a[1]~q ;
wire \add_in_r_b[0]~q ;
wire \Add1~2_combout ;
wire \add_in_r_a[0]~q ;
wire \add_in_r_d[9]~q ;
wire \Add3~3_combout ;
wire \add_in_r_c[9]~q ;
wire \add_in_r_d[8]~q ;
wire \Add3~4_combout ;
wire \add_in_r_c[8]~q ;
wire \add_in_r_d[7]~q ;
wire \Add3~5_combout ;
wire \add_in_r_c[7]~q ;
wire \add_in_r_d[6]~q ;
wire \Add3~6_combout ;
wire \add_in_r_c[6]~q ;
wire \add_in_r_d[5]~q ;
wire \Add3~7_combout ;
wire \add_in_r_c[5]~q ;
wire \add_in_r_d[4]~q ;
wire \Add3~8_combout ;
wire \add_in_r_c[4]~q ;
wire \add_in_r_d[3]~q ;
wire \Add3~9_combout ;
wire \add_in_r_c[3]~q ;
wire \add_in_r_b[9]~q ;
wire \Add1~3_combout ;
wire \add_in_r_a[9]~q ;
wire \add_in_r_b[8]~q ;
wire \Add1~4_combout ;
wire \add_in_r_a[8]~q ;
wire \add_in_r_b[7]~q ;
wire \Add1~5_combout ;
wire \add_in_r_a[7]~q ;
wire \add_in_r_b[6]~q ;
wire \Add1~6_combout ;
wire \add_in_r_a[6]~q ;
wire \add_in_r_b[5]~q ;
wire \Add1~7_combout ;
wire \add_in_r_a[5]~q ;
wire \add_in_r_b[4]~q ;
wire \Add1~8_combout ;
wire \add_in_r_a[4]~q ;
wire \add_in_r_b[3]~q ;
wire \Add1~9_combout ;
wire \add_in_r_a[3]~q ;
wire \sign_sel[0]~q ;
wire \sign_sel[1]~q ;
wire \Mux0~0_combout ;
wire \add_in_i_d~0_combout ;
wire \add_in_i_c~0_combout ;
wire \add_in_i_d~1_combout ;
wire \add_in_i_c~1_combout ;
wire \add_in_i_d~2_combout ;
wire \add_in_i_c~2_combout ;
wire \add_in_i_d~3_combout ;
wire \add_in_i_c~3_combout ;
wire \add_in_i_d~4_combout ;
wire \add_in_i_c~4_combout ;
wire \add_in_i_d~5_combout ;
wire \add_in_i_c~5_combout ;
wire \add_in_i_d~6_combout ;
wire \add_in_i_c~6_combout ;
wire \add_in_i_d~7_combout ;
wire \add_in_i_c~7_combout ;
wire \add_in_i_d~8_combout ;
wire \add_in_i_c~8_combout ;
wire \add_in_i_d~9_combout ;
wire \add_in_i_c~9_combout ;
wire \add_in_r_d~0_combout ;
wire \add_in_r_c~0_combout ;
wire \add_in_r_d~1_combout ;
wire \add_in_r_c~1_combout ;
wire \add_in_r_d~2_combout ;
wire \add_in_r_c~2_combout ;
wire \add_in_r_d~3_combout ;
wire \add_in_r_c~3_combout ;
wire \add_in_r_d~4_combout ;
wire \add_in_r_c~4_combout ;
wire \add_in_r_d~5_combout ;
wire \add_in_r_c~5_combout ;
wire \add_in_r_d~6_combout ;
wire \add_in_r_c~6_combout ;
wire \add_in_r_d~7_combout ;
wire \add_in_r_c~7_combout ;
wire \add_in_r_d~8_combout ;
wire \add_in_r_c~8_combout ;
wire \add_in_r_d~9_combout ;
wire \add_in_r_c~9_combout ;
wire \offset_counter[5]~28_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \data_val_i~0_combout ;
wire \sign_vec[3]~1_combout ;
wire \sign_vec[1]~2_combout ;
wire \data_real_o~0_combout ;
wire \data_real_o~1_combout ;
wire \data_real_o~2_combout ;
wire \data_real_o~3_combout ;
wire \data_real_o~4_combout ;
wire \data_real_o~5_combout ;
wire \data_real_o~6_combout ;
wire \data_real_o~7_combout ;
wire \data_real_o~8_combout ;
wire \data_real_o~9_combout ;


fftsign_asj_fft_pround_15 \gen_full_rnd:u1 (
	.pipeline_dffe_2(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.output_i_2(\output_i[2]~q ),
	.output_i_1(\output_i[1]~q ),
	.output_i_0(\output_i[0]~q ),
	.output_i_11(\output_i[11]~q ),
	.output_i_3(\output_i[3]~q ),
	.output_i_4(\output_i[4]~q ),
	.output_i_5(\output_i[5]~q ),
	.output_i_6(\output_i[6]~q ),
	.output_i_7(\output_i[7]~q ),
	.output_i_8(\output_i[8]~q ),
	.output_i_9(\output_i[9]~q ),
	.output_i_10(\output_i[10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_pround_14 \gen_full_rnd:u0 (
	.pipeline_dffe_2(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.output_r_2(\output_r[2]~q ),
	.output_r_1(\output_r[1]~q ),
	.output_r_0(\output_r[0]~q ),
	.output_r_11(\output_r[11]~q ),
	.output_r_3(\output_r[3]~q ),
	.output_r_4(\output_r[4]~q ),
	.output_r_5(\output_r[5]~q ),
	.output_r_6(\output_r[6]~q ),
	.output_r_7(\output_r[7]~q ),
	.output_r_8(\output_r[8]~q ),
	.output_r_9(\output_r[9]~q ),
	.output_r_10(\output_r[10]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

fftsign_asj_fft_tdl_bit_1 \gen_burst_val:delay_val (
	.data_in(\data_val_i~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_4(tdl_arr_41),
	.clk(clk));

dffeas \output_i[2] (
	.clk(clk),
	.d(\output_i[2]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[2]~q ),
	.prn(vcc));
defparam \output_i[2] .is_wysiwyg = "true";
defparam \output_i[2] .power_up = "low";

dffeas \output_i[1] (
	.clk(clk),
	.d(\output_i[1]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[1]~q ),
	.prn(vcc));
defparam \output_i[1] .is_wysiwyg = "true";
defparam \output_i[1] .power_up = "low";

dffeas \output_i[0] (
	.clk(clk),
	.d(\output_i[0]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[0]~q ),
	.prn(vcc));
defparam \output_i[0] .is_wysiwyg = "true";
defparam \output_i[0] .power_up = "low";

dffeas \output_i[11] (
	.clk(clk),
	.d(\output_i[11]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[11]~q ),
	.prn(vcc));
defparam \output_i[11] .is_wysiwyg = "true";
defparam \output_i[11] .power_up = "low";

dffeas \output_r[2] (
	.clk(clk),
	.d(\output_r[2]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[2]~q ),
	.prn(vcc));
defparam \output_r[2] .is_wysiwyg = "true";
defparam \output_r[2] .power_up = "low";

dffeas \output_r[1] (
	.clk(clk),
	.d(\output_r[1]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[1]~q ),
	.prn(vcc));
defparam \output_r[1] .is_wysiwyg = "true";
defparam \output_r[1] .power_up = "low";

dffeas \output_r[0] (
	.clk(clk),
	.d(\output_r[0]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[0]~q ),
	.prn(vcc));
defparam \output_r[0] .is_wysiwyg = "true";
defparam \output_r[0] .power_up = "low";

dffeas \output_r[11] (
	.clk(clk),
	.d(\output_r[11]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[11]~q ),
	.prn(vcc));
defparam \output_r[11] .is_wysiwyg = "true";
defparam \output_r[11] .power_up = "low";

dffeas \output_i[3] (
	.clk(clk),
	.d(\output_i[3]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[3]~q ),
	.prn(vcc));
defparam \output_i[3] .is_wysiwyg = "true";
defparam \output_i[3] .power_up = "low";

dffeas \output_r[3] (
	.clk(clk),
	.d(\output_r[3]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[3]~q ),
	.prn(vcc));
defparam \output_r[3] .is_wysiwyg = "true";
defparam \output_r[3] .power_up = "low";

dffeas \output_i[4] (
	.clk(clk),
	.d(\output_i[4]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[4]~q ),
	.prn(vcc));
defparam \output_i[4] .is_wysiwyg = "true";
defparam \output_i[4] .power_up = "low";

dffeas \output_r[4] (
	.clk(clk),
	.d(\output_r[4]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[4]~q ),
	.prn(vcc));
defparam \output_r[4] .is_wysiwyg = "true";
defparam \output_r[4] .power_up = "low";

dffeas \output_i[5] (
	.clk(clk),
	.d(\output_i[5]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[5]~q ),
	.prn(vcc));
defparam \output_i[5] .is_wysiwyg = "true";
defparam \output_i[5] .power_up = "low";

dffeas \output_r[5] (
	.clk(clk),
	.d(\output_r[5]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[5]~q ),
	.prn(vcc));
defparam \output_r[5] .is_wysiwyg = "true";
defparam \output_r[5] .power_up = "low";

dffeas \output_i[6] (
	.clk(clk),
	.d(\output_i[6]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[6]~q ),
	.prn(vcc));
defparam \output_i[6] .is_wysiwyg = "true";
defparam \output_i[6] .power_up = "low";

dffeas \output_r[6] (
	.clk(clk),
	.d(\output_r[6]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[6]~q ),
	.prn(vcc));
defparam \output_r[6] .is_wysiwyg = "true";
defparam \output_r[6] .power_up = "low";

dffeas \output_i[7] (
	.clk(clk),
	.d(\output_i[7]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[7]~q ),
	.prn(vcc));
defparam \output_i[7] .is_wysiwyg = "true";
defparam \output_i[7] .power_up = "low";

dffeas \output_r[7] (
	.clk(clk),
	.d(\output_r[7]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[7]~q ),
	.prn(vcc));
defparam \output_r[7] .is_wysiwyg = "true";
defparam \output_r[7] .power_up = "low";

dffeas \output_i[8] (
	.clk(clk),
	.d(\output_i[8]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[8]~q ),
	.prn(vcc));
defparam \output_i[8] .is_wysiwyg = "true";
defparam \output_i[8] .power_up = "low";

dffeas \output_r[8] (
	.clk(clk),
	.d(\output_r[8]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[8]~q ),
	.prn(vcc));
defparam \output_r[8] .is_wysiwyg = "true";
defparam \output_r[8] .power_up = "low";

dffeas \output_i[9] (
	.clk(clk),
	.d(\output_i[9]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[9]~q ),
	.prn(vcc));
defparam \output_i[9] .is_wysiwyg = "true";
defparam \output_i[9] .power_up = "low";

dffeas \output_r[9] (
	.clk(clk),
	.d(\output_r[9]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[9]~q ),
	.prn(vcc));
defparam \output_r[9] .is_wysiwyg = "true";
defparam \output_r[9] .power_up = "low";

dffeas \output_i[10] (
	.clk(clk),
	.d(\output_i[10]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_i[10]~q ),
	.prn(vcc));
defparam \output_i[10] .is_wysiwyg = "true";
defparam \output_i[10] .power_up = "low";

dffeas \output_r[10] (
	.clk(clk),
	.d(\output_r[10]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\output_r[10]~q ),
	.prn(vcc));
defparam \output_r[10] .is_wysiwyg = "true";
defparam \output_r[10] .power_up = "low";

dffeas \result_ib[2] (
	.clk(clk),
	.d(\result_ib[2]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[2]~q ),
	.prn(vcc));
defparam \result_ib[2] .is_wysiwyg = "true";
defparam \result_ib[2] .power_up = "low";

dffeas \result_ia[2] (
	.clk(clk),
	.d(\result_ia[2]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[2]~q ),
	.prn(vcc));
defparam \result_ia[2] .is_wysiwyg = "true";
defparam \result_ia[2] .power_up = "low";

dffeas \result_ib[1] (
	.clk(clk),
	.d(\result_ib[1]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[1]~q ),
	.prn(vcc));
defparam \result_ib[1] .is_wysiwyg = "true";
defparam \result_ib[1] .power_up = "low";

dffeas \result_ia[1] (
	.clk(clk),
	.d(\result_ia[1]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[1]~q ),
	.prn(vcc));
defparam \result_ia[1] .is_wysiwyg = "true";
defparam \result_ia[1] .power_up = "low";

dffeas \result_ib[0] (
	.clk(clk),
	.d(\result_ib[0]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[0]~q ),
	.prn(vcc));
defparam \result_ib[0] .is_wysiwyg = "true";
defparam \result_ib[0] .power_up = "low";

dffeas \result_ia[0] (
	.clk(clk),
	.d(\result_ia[0]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[0]~q ),
	.prn(vcc));
defparam \result_ia[0] .is_wysiwyg = "true";
defparam \result_ia[0] .power_up = "low";

cycloneive_lcell_comb \output_i[0]~13 (
	.dataa(\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\output_i[0]~13_cout ));
defparam \output_i[0]~13 .lut_mask = 16'h0055;
defparam \output_i[0]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \output_i[0]~14 (
	.dataa(\Add11~2_combout ),
	.datab(\result_ia[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[0]~13_cout ),
	.combout(\output_i[0]~14_combout ),
	.cout(\output_i[0]~15 ));
defparam \output_i[0]~14 .lut_mask = 16'h96BF;
defparam \output_i[0]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[1]~16 (
	.dataa(\Add11~1_combout ),
	.datab(\result_ia[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[0]~15 ),
	.combout(\output_i[1]~16_combout ),
	.cout(\output_i[1]~17 ));
defparam \output_i[1]~16 .lut_mask = 16'h96DF;
defparam \output_i[1]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[2]~18 (
	.dataa(\Add11~0_combout ),
	.datab(\result_ia[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[1]~17 ),
	.combout(\output_i[2]~18_combout ),
	.cout(\output_i[2]~19 ));
defparam \output_i[2]~18 .lut_mask = 16'h96BF;
defparam \output_i[2]~18 .sum_lutc_input = "cin";

dffeas \result_ib[10] (
	.clk(clk),
	.d(\result_ib[10]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[10]~q ),
	.prn(vcc));
defparam \result_ib[10] .is_wysiwyg = "true";
defparam \result_ib[10] .power_up = "low";

dffeas \result_ia[10] (
	.clk(clk),
	.d(\result_ia[10]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[10]~q ),
	.prn(vcc));
defparam \result_ia[10] .is_wysiwyg = "true";
defparam \result_ia[10] .power_up = "low";

dffeas \result_ib[9] (
	.clk(clk),
	.d(\result_ib[9]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[9]~q ),
	.prn(vcc));
defparam \result_ib[9] .is_wysiwyg = "true";
defparam \result_ib[9] .power_up = "low";

dffeas \result_ia[9] (
	.clk(clk),
	.d(\result_ia[9]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[9]~q ),
	.prn(vcc));
defparam \result_ia[9] .is_wysiwyg = "true";
defparam \result_ia[9] .power_up = "low";

dffeas \result_ib[8] (
	.clk(clk),
	.d(\result_ib[8]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[8]~q ),
	.prn(vcc));
defparam \result_ib[8] .is_wysiwyg = "true";
defparam \result_ib[8] .power_up = "low";

dffeas \result_ia[8] (
	.clk(clk),
	.d(\result_ia[8]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[8]~q ),
	.prn(vcc));
defparam \result_ia[8] .is_wysiwyg = "true";
defparam \result_ia[8] .power_up = "low";

dffeas \result_ib[7] (
	.clk(clk),
	.d(\result_ib[7]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[7]~q ),
	.prn(vcc));
defparam \result_ib[7] .is_wysiwyg = "true";
defparam \result_ib[7] .power_up = "low";

dffeas \result_ia[7] (
	.clk(clk),
	.d(\result_ia[7]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[7]~q ),
	.prn(vcc));
defparam \result_ia[7] .is_wysiwyg = "true";
defparam \result_ia[7] .power_up = "low";

dffeas \result_ib[6] (
	.clk(clk),
	.d(\result_ib[6]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[6]~q ),
	.prn(vcc));
defparam \result_ib[6] .is_wysiwyg = "true";
defparam \result_ib[6] .power_up = "low";

dffeas \result_ia[6] (
	.clk(clk),
	.d(\result_ia[6]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[6]~q ),
	.prn(vcc));
defparam \result_ia[6] .is_wysiwyg = "true";
defparam \result_ia[6] .power_up = "low";

dffeas \result_ib[5] (
	.clk(clk),
	.d(\result_ib[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[5]~q ),
	.prn(vcc));
defparam \result_ib[5] .is_wysiwyg = "true";
defparam \result_ib[5] .power_up = "low";

dffeas \result_ia[5] (
	.clk(clk),
	.d(\result_ia[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[5]~q ),
	.prn(vcc));
defparam \result_ia[5] .is_wysiwyg = "true";
defparam \result_ia[5] .power_up = "low";

dffeas \result_ib[4] (
	.clk(clk),
	.d(\result_ib[4]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[4]~q ),
	.prn(vcc));
defparam \result_ib[4] .is_wysiwyg = "true";
defparam \result_ib[4] .power_up = "low";

dffeas \result_ia[4] (
	.clk(clk),
	.d(\result_ia[4]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[4]~q ),
	.prn(vcc));
defparam \result_ia[4] .is_wysiwyg = "true";
defparam \result_ia[4] .power_up = "low";

dffeas \result_ib[3] (
	.clk(clk),
	.d(\result_ib[3]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ib[3]~q ),
	.prn(vcc));
defparam \result_ib[3] .is_wysiwyg = "true";
defparam \result_ib[3] .power_up = "low";

dffeas \result_ia[3] (
	.clk(clk),
	.d(\result_ia[3]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ia[3]~q ),
	.prn(vcc));
defparam \result_ia[3] .is_wysiwyg = "true";
defparam \result_ia[3] .power_up = "low";

cycloneive_lcell_comb \output_i[3]~20 (
	.dataa(\Add11~10_combout ),
	.datab(\result_ia[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[2]~19 ),
	.combout(\output_i[3]~20_combout ),
	.cout(\output_i[3]~21 ));
defparam \output_i[3]~20 .lut_mask = 16'h96DF;
defparam \output_i[3]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[4]~22 (
	.dataa(\Add11~9_combout ),
	.datab(\result_ia[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[3]~21 ),
	.combout(\output_i[4]~22_combout ),
	.cout(\output_i[4]~23 ));
defparam \output_i[4]~22 .lut_mask = 16'h96BF;
defparam \output_i[4]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[5]~24 (
	.dataa(\Add11~8_combout ),
	.datab(\result_ia[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[4]~23 ),
	.combout(\output_i[5]~24_combout ),
	.cout(\output_i[5]~25 ));
defparam \output_i[5]~24 .lut_mask = 16'h96DF;
defparam \output_i[5]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[6]~26 (
	.dataa(\Add11~7_combout ),
	.datab(\result_ia[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[5]~25 ),
	.combout(\output_i[6]~26_combout ),
	.cout(\output_i[6]~27 ));
defparam \output_i[6]~26 .lut_mask = 16'h96BF;
defparam \output_i[6]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[7]~28 (
	.dataa(\Add11~6_combout ),
	.datab(\result_ia[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[6]~27 ),
	.combout(\output_i[7]~28_combout ),
	.cout(\output_i[7]~29 ));
defparam \output_i[7]~28 .lut_mask = 16'h96DF;
defparam \output_i[7]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[8]~30 (
	.dataa(\Add11~5_combout ),
	.datab(\result_ia[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[7]~29 ),
	.combout(\output_i[8]~30_combout ),
	.cout(\output_i[8]~31 ));
defparam \output_i[8]~30 .lut_mask = 16'h96BF;
defparam \output_i[8]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[9]~32 (
	.dataa(\Add11~4_combout ),
	.datab(\result_ia[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[8]~31 ),
	.combout(\output_i[9]~32_combout ),
	.cout(\output_i[9]~33 ));
defparam \output_i[9]~32 .lut_mask = 16'h96DF;
defparam \output_i[9]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[10]~34 (
	.dataa(\Add11~3_combout ),
	.datab(\result_ia[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_i[9]~33 ),
	.combout(\output_i[10]~34_combout ),
	.cout(\output_i[10]~35 ));
defparam \output_i[10]~34 .lut_mask = 16'h96BF;
defparam \output_i[10]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_i[11]~36 (
	.dataa(\Add11~3_combout ),
	.datab(\result_ia[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\output_i[10]~35 ),
	.combout(\output_i[11]~36_combout ),
	.cout());
defparam \output_i[11]~36 .lut_mask = 16'h9696;
defparam \output_i[11]~36 .sum_lutc_input = "cin";

dffeas \result_rb[2] (
	.clk(clk),
	.d(\result_rb[2]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[2]~q ),
	.prn(vcc));
defparam \result_rb[2] .is_wysiwyg = "true";
defparam \result_rb[2] .power_up = "low";

dffeas \result_ra[2] (
	.clk(clk),
	.d(\result_ra[2]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[2]~q ),
	.prn(vcc));
defparam \result_ra[2] .is_wysiwyg = "true";
defparam \result_ra[2] .power_up = "low";

dffeas \result_rb[1] (
	.clk(clk),
	.d(\result_rb[1]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[1]~q ),
	.prn(vcc));
defparam \result_rb[1] .is_wysiwyg = "true";
defparam \result_rb[1] .power_up = "low";

dffeas \result_ra[1] (
	.clk(clk),
	.d(\result_ra[1]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[1]~q ),
	.prn(vcc));
defparam \result_ra[1] .is_wysiwyg = "true";
defparam \result_ra[1] .power_up = "low";

dffeas \result_rb[0] (
	.clk(clk),
	.d(\result_rb[0]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[0]~q ),
	.prn(vcc));
defparam \result_rb[0] .is_wysiwyg = "true";
defparam \result_rb[0] .power_up = "low";

dffeas \result_ra[0] (
	.clk(clk),
	.d(\result_ra[0]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[0]~q ),
	.prn(vcc));
defparam \result_ra[0] .is_wysiwyg = "true";
defparam \result_ra[0] .power_up = "low";

cycloneive_lcell_comb \output_r[0]~13 (
	.dataa(\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\output_r[0]~13_cout ));
defparam \output_r[0]~13 .lut_mask = 16'h0055;
defparam \output_r[0]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \output_r[0]~14 (
	.dataa(\Add9~2_combout ),
	.datab(\result_ra[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[0]~13_cout ),
	.combout(\output_r[0]~14_combout ),
	.cout(\output_r[0]~15 ));
defparam \output_r[0]~14 .lut_mask = 16'h96BF;
defparam \output_r[0]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[1]~16 (
	.dataa(\Add9~1_combout ),
	.datab(\result_ra[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[0]~15 ),
	.combout(\output_r[1]~16_combout ),
	.cout(\output_r[1]~17 ));
defparam \output_r[1]~16 .lut_mask = 16'h96DF;
defparam \output_r[1]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[2]~18 (
	.dataa(\Add9~0_combout ),
	.datab(\result_ra[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[1]~17 ),
	.combout(\output_r[2]~18_combout ),
	.cout(\output_r[2]~19 ));
defparam \output_r[2]~18 .lut_mask = 16'h96BF;
defparam \output_r[2]~18 .sum_lutc_input = "cin";

dffeas \result_rb[10] (
	.clk(clk),
	.d(\result_rb[10]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[10]~q ),
	.prn(vcc));
defparam \result_rb[10] .is_wysiwyg = "true";
defparam \result_rb[10] .power_up = "low";

dffeas \result_ra[10] (
	.clk(clk),
	.d(\result_ra[10]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[10]~q ),
	.prn(vcc));
defparam \result_ra[10] .is_wysiwyg = "true";
defparam \result_ra[10] .power_up = "low";

dffeas \result_rb[9] (
	.clk(clk),
	.d(\result_rb[9]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[9]~q ),
	.prn(vcc));
defparam \result_rb[9] .is_wysiwyg = "true";
defparam \result_rb[9] .power_up = "low";

dffeas \result_ra[9] (
	.clk(clk),
	.d(\result_ra[9]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[9]~q ),
	.prn(vcc));
defparam \result_ra[9] .is_wysiwyg = "true";
defparam \result_ra[9] .power_up = "low";

dffeas \result_rb[8] (
	.clk(clk),
	.d(\result_rb[8]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[8]~q ),
	.prn(vcc));
defparam \result_rb[8] .is_wysiwyg = "true";
defparam \result_rb[8] .power_up = "low";

dffeas \result_ra[8] (
	.clk(clk),
	.d(\result_ra[8]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[8]~q ),
	.prn(vcc));
defparam \result_ra[8] .is_wysiwyg = "true";
defparam \result_ra[8] .power_up = "low";

dffeas \result_rb[7] (
	.clk(clk),
	.d(\result_rb[7]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[7]~q ),
	.prn(vcc));
defparam \result_rb[7] .is_wysiwyg = "true";
defparam \result_rb[7] .power_up = "low";

dffeas \result_ra[7] (
	.clk(clk),
	.d(\result_ra[7]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[7]~q ),
	.prn(vcc));
defparam \result_ra[7] .is_wysiwyg = "true";
defparam \result_ra[7] .power_up = "low";

dffeas \result_rb[6] (
	.clk(clk),
	.d(\result_rb[6]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[6]~q ),
	.prn(vcc));
defparam \result_rb[6] .is_wysiwyg = "true";
defparam \result_rb[6] .power_up = "low";

dffeas \result_ra[6] (
	.clk(clk),
	.d(\result_ra[6]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[6]~q ),
	.prn(vcc));
defparam \result_ra[6] .is_wysiwyg = "true";
defparam \result_ra[6] .power_up = "low";

dffeas \result_rb[5] (
	.clk(clk),
	.d(\result_rb[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[5]~q ),
	.prn(vcc));
defparam \result_rb[5] .is_wysiwyg = "true";
defparam \result_rb[5] .power_up = "low";

dffeas \result_ra[5] (
	.clk(clk),
	.d(\result_ra[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[5]~q ),
	.prn(vcc));
defparam \result_ra[5] .is_wysiwyg = "true";
defparam \result_ra[5] .power_up = "low";

dffeas \result_rb[4] (
	.clk(clk),
	.d(\result_rb[4]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[4]~q ),
	.prn(vcc));
defparam \result_rb[4] .is_wysiwyg = "true";
defparam \result_rb[4] .power_up = "low";

dffeas \result_ra[4] (
	.clk(clk),
	.d(\result_ra[4]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[4]~q ),
	.prn(vcc));
defparam \result_ra[4] .is_wysiwyg = "true";
defparam \result_ra[4] .power_up = "low";

dffeas \result_rb[3] (
	.clk(clk),
	.d(\result_rb[3]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_rb[3]~q ),
	.prn(vcc));
defparam \result_rb[3] .is_wysiwyg = "true";
defparam \result_rb[3] .power_up = "low";

dffeas \result_ra[3] (
	.clk(clk),
	.d(\result_ra[3]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\result_ra[3]~q ),
	.prn(vcc));
defparam \result_ra[3] .is_wysiwyg = "true";
defparam \result_ra[3] .power_up = "low";

cycloneive_lcell_comb \output_r[3]~20 (
	.dataa(\Add9~10_combout ),
	.datab(\result_ra[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[2]~19 ),
	.combout(\output_r[3]~20_combout ),
	.cout(\output_r[3]~21 ));
defparam \output_r[3]~20 .lut_mask = 16'h96DF;
defparam \output_r[3]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[4]~22 (
	.dataa(\Add9~9_combout ),
	.datab(\result_ra[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[3]~21 ),
	.combout(\output_r[4]~22_combout ),
	.cout(\output_r[4]~23 ));
defparam \output_r[4]~22 .lut_mask = 16'h96BF;
defparam \output_r[4]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[5]~24 (
	.dataa(\Add9~8_combout ),
	.datab(\result_ra[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[4]~23 ),
	.combout(\output_r[5]~24_combout ),
	.cout(\output_r[5]~25 ));
defparam \output_r[5]~24 .lut_mask = 16'h96DF;
defparam \output_r[5]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[6]~26 (
	.dataa(\Add9~7_combout ),
	.datab(\result_ra[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[5]~25 ),
	.combout(\output_r[6]~26_combout ),
	.cout(\output_r[6]~27 ));
defparam \output_r[6]~26 .lut_mask = 16'h96BF;
defparam \output_r[6]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[7]~28 (
	.dataa(\Add9~6_combout ),
	.datab(\result_ra[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[6]~27 ),
	.combout(\output_r[7]~28_combout ),
	.cout(\output_r[7]~29 ));
defparam \output_r[7]~28 .lut_mask = 16'h96DF;
defparam \output_r[7]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[8]~30 (
	.dataa(\Add9~5_combout ),
	.datab(\result_ra[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[7]~29 ),
	.combout(\output_r[8]~30_combout ),
	.cout(\output_r[8]~31 ));
defparam \output_r[8]~30 .lut_mask = 16'h96BF;
defparam \output_r[8]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[9]~32 (
	.dataa(\Add9~4_combout ),
	.datab(\result_ra[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[8]~31 ),
	.combout(\output_r[9]~32_combout ),
	.cout(\output_r[9]~33 ));
defparam \output_r[9]~32 .lut_mask = 16'h96DF;
defparam \output_r[9]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[10]~34 (
	.dataa(\Add9~3_combout ),
	.datab(\result_ra[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\output_r[9]~33 ),
	.combout(\output_r[10]~34_combout ),
	.cout(\output_r[10]~35 ));
defparam \output_r[10]~34 .lut_mask = 16'h96BF;
defparam \output_r[10]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \output_r[11]~36 (
	.dataa(\Add9~3_combout ),
	.datab(\result_ra[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\output_r[10]~35 ),
	.combout(\output_r[11]~36_combout ),
	.cout());
defparam \output_r[11]~36 .lut_mask = 16'h9696;
defparam \output_r[11]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[0]~12 (
	.dataa(\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_ib[0]~12_cout ));
defparam \result_ib[0]~12 .lut_mask = 16'h0055;
defparam \result_ib[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_ib[0]~13 (
	.dataa(\Add4~2_combout ),
	.datab(\add_in_i_c[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[0]~12_cout ),
	.combout(\result_ib[0]~13_combout ),
	.cout(\result_ib[0]~14 ));
defparam \result_ib[0]~13 .lut_mask = 16'h96BF;
defparam \result_ib[0]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[1]~15 (
	.dataa(\Add4~1_combout ),
	.datab(\add_in_i_c[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[0]~14 ),
	.combout(\result_ib[1]~15_combout ),
	.cout(\result_ib[1]~16 ));
defparam \result_ib[1]~15 .lut_mask = 16'h96DF;
defparam \result_ib[1]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[2]~17 (
	.dataa(\Add4~0_combout ),
	.datab(\add_in_i_c[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[1]~16 ),
	.combout(\result_ib[2]~17_combout ),
	.cout(\result_ib[2]~18 ));
defparam \result_ib[2]~17 .lut_mask = 16'h96BF;
defparam \result_ib[2]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[0]~12 (
	.dataa(\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_ia[0]~12_cout ));
defparam \result_ia[0]~12 .lut_mask = 16'h0055;
defparam \result_ia[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_ia[0]~13 (
	.dataa(\Add2~2_combout ),
	.datab(\add_in_i_a[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[0]~12_cout ),
	.combout(\result_ia[0]~13_combout ),
	.cout(\result_ia[0]~14 ));
defparam \result_ia[0]~13 .lut_mask = 16'h96BF;
defparam \result_ia[0]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[1]~15 (
	.dataa(\Add2~1_combout ),
	.datab(\add_in_i_a[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[0]~14 ),
	.combout(\result_ia[1]~15_combout ),
	.cout(\result_ia[1]~16 ));
defparam \result_ia[1]~15 .lut_mask = 16'h96DF;
defparam \result_ia[1]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[2]~17 (
	.dataa(\Add2~0_combout ),
	.datab(\add_in_i_a[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[1]~16 ),
	.combout(\result_ia[2]~17_combout ),
	.cout(\result_ia[2]~18 ));
defparam \result_ia[2]~17 .lut_mask = 16'h96BF;
defparam \result_ia[2]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[3]~19 (
	.dataa(\Add4~9_combout ),
	.datab(\add_in_i_c[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[2]~18 ),
	.combout(\result_ib[3]~19_combout ),
	.cout(\result_ib[3]~20 ));
defparam \result_ib[3]~19 .lut_mask = 16'h96DF;
defparam \result_ib[3]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[4]~21 (
	.dataa(\Add4~8_combout ),
	.datab(\add_in_i_c[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[3]~20 ),
	.combout(\result_ib[4]~21_combout ),
	.cout(\result_ib[4]~22 ));
defparam \result_ib[4]~21 .lut_mask = 16'h96BF;
defparam \result_ib[4]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[5]~23 (
	.dataa(\Add4~7_combout ),
	.datab(\add_in_i_c[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[4]~22 ),
	.combout(\result_ib[5]~23_combout ),
	.cout(\result_ib[5]~24 ));
defparam \result_ib[5]~23 .lut_mask = 16'h96DF;
defparam \result_ib[5]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[6]~25 (
	.dataa(\Add4~6_combout ),
	.datab(\add_in_i_c[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[5]~24 ),
	.combout(\result_ib[6]~25_combout ),
	.cout(\result_ib[6]~26 ));
defparam \result_ib[6]~25 .lut_mask = 16'h96BF;
defparam \result_ib[6]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[7]~27 (
	.dataa(\Add4~5_combout ),
	.datab(\add_in_i_c[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[6]~26 ),
	.combout(\result_ib[7]~27_combout ),
	.cout(\result_ib[7]~28 ));
defparam \result_ib[7]~27 .lut_mask = 16'h96DF;
defparam \result_ib[7]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[8]~29 (
	.dataa(\Add4~4_combout ),
	.datab(\add_in_i_c[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[7]~28 ),
	.combout(\result_ib[8]~29_combout ),
	.cout(\result_ib[8]~30 ));
defparam \result_ib[8]~29 .lut_mask = 16'h96BF;
defparam \result_ib[8]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[9]~31 (
	.dataa(\Add4~3_combout ),
	.datab(\add_in_i_c[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ib[8]~30 ),
	.combout(\result_ib[9]~31_combout ),
	.cout(\result_ib[9]~32 ));
defparam \result_ib[9]~31 .lut_mask = 16'h96DF;
defparam \result_ib[9]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ib[10]~33 (
	.dataa(\Add4~3_combout ),
	.datab(\add_in_i_c[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_ib[9]~32 ),
	.combout(\result_ib[10]~33_combout ),
	.cout());
defparam \result_ib[10]~33 .lut_mask = 16'h9696;
defparam \result_ib[10]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[3]~19 (
	.dataa(\Add2~9_combout ),
	.datab(\add_in_i_a[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[2]~18 ),
	.combout(\result_ia[3]~19_combout ),
	.cout(\result_ia[3]~20 ));
defparam \result_ia[3]~19 .lut_mask = 16'h96DF;
defparam \result_ia[3]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[4]~21 (
	.dataa(\Add2~8_combout ),
	.datab(\add_in_i_a[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[3]~20 ),
	.combout(\result_ia[4]~21_combout ),
	.cout(\result_ia[4]~22 ));
defparam \result_ia[4]~21 .lut_mask = 16'h96BF;
defparam \result_ia[4]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[5]~23 (
	.dataa(\Add2~7_combout ),
	.datab(\add_in_i_a[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[4]~22 ),
	.combout(\result_ia[5]~23_combout ),
	.cout(\result_ia[5]~24 ));
defparam \result_ia[5]~23 .lut_mask = 16'h96DF;
defparam \result_ia[5]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[6]~25 (
	.dataa(\Add2~6_combout ),
	.datab(\add_in_i_a[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[5]~24 ),
	.combout(\result_ia[6]~25_combout ),
	.cout(\result_ia[6]~26 ));
defparam \result_ia[6]~25 .lut_mask = 16'h96BF;
defparam \result_ia[6]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[7]~27 (
	.dataa(\Add2~5_combout ),
	.datab(\add_in_i_a[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[6]~26 ),
	.combout(\result_ia[7]~27_combout ),
	.cout(\result_ia[7]~28 ));
defparam \result_ia[7]~27 .lut_mask = 16'h96DF;
defparam \result_ia[7]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[8]~29 (
	.dataa(\Add2~4_combout ),
	.datab(\add_in_i_a[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[7]~28 ),
	.combout(\result_ia[8]~29_combout ),
	.cout(\result_ia[8]~30 ));
defparam \result_ia[8]~29 .lut_mask = 16'h96BF;
defparam \result_ia[8]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[9]~31 (
	.dataa(\Add2~3_combout ),
	.datab(\add_in_i_a[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ia[8]~30 ),
	.combout(\result_ia[9]~31_combout ),
	.cout(\result_ia[9]~32 ));
defparam \result_ia[9]~31 .lut_mask = 16'h96DF;
defparam \result_ia[9]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ia[10]~33 (
	.dataa(\Add2~3_combout ),
	.datab(\add_in_i_a[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_ia[9]~32 ),
	.combout(\result_ia[10]~33_combout ),
	.cout());
defparam \result_ia[10]~33 .lut_mask = 16'h9696;
defparam \result_ia[10]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[0]~12 (
	.dataa(\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_rb[0]~12_cout ));
defparam \result_rb[0]~12 .lut_mask = 16'h0055;
defparam \result_rb[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_rb[0]~13 (
	.dataa(\Add3~2_combout ),
	.datab(\add_in_r_c[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[0]~12_cout ),
	.combout(\result_rb[0]~13_combout ),
	.cout(\result_rb[0]~14 ));
defparam \result_rb[0]~13 .lut_mask = 16'h96BF;
defparam \result_rb[0]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[1]~15 (
	.dataa(\Add3~1_combout ),
	.datab(\add_in_r_c[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[0]~14 ),
	.combout(\result_rb[1]~15_combout ),
	.cout(\result_rb[1]~16 ));
defparam \result_rb[1]~15 .lut_mask = 16'h96DF;
defparam \result_rb[1]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[2]~17 (
	.dataa(\Add3~0_combout ),
	.datab(\add_in_r_c[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[1]~16 ),
	.combout(\result_rb[2]~17_combout ),
	.cout(\result_rb[2]~18 ));
defparam \result_rb[2]~17 .lut_mask = 16'h96BF;
defparam \result_rb[2]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[0]~12 (
	.dataa(\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\result_ra[0]~12_cout ));
defparam \result_ra[0]~12 .lut_mask = 16'h0055;
defparam \result_ra[0]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \result_ra[0]~13 (
	.dataa(\Add1~2_combout ),
	.datab(\add_in_r_a[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[0]~12_cout ),
	.combout(\result_ra[0]~13_combout ),
	.cout(\result_ra[0]~14 ));
defparam \result_ra[0]~13 .lut_mask = 16'h96BF;
defparam \result_ra[0]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[1]~15 (
	.dataa(\Add1~1_combout ),
	.datab(\add_in_r_a[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[0]~14 ),
	.combout(\result_ra[1]~15_combout ),
	.cout(\result_ra[1]~16 ));
defparam \result_ra[1]~15 .lut_mask = 16'h96DF;
defparam \result_ra[1]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[2]~17 (
	.dataa(\Add1~0_combout ),
	.datab(\add_in_r_a[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[1]~16 ),
	.combout(\result_ra[2]~17_combout ),
	.cout(\result_ra[2]~18 ));
defparam \result_ra[2]~17 .lut_mask = 16'h96BF;
defparam \result_ra[2]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[3]~19 (
	.dataa(\Add3~9_combout ),
	.datab(\add_in_r_c[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[2]~18 ),
	.combout(\result_rb[3]~19_combout ),
	.cout(\result_rb[3]~20 ));
defparam \result_rb[3]~19 .lut_mask = 16'h96DF;
defparam \result_rb[3]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[4]~21 (
	.dataa(\Add3~8_combout ),
	.datab(\add_in_r_c[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[3]~20 ),
	.combout(\result_rb[4]~21_combout ),
	.cout(\result_rb[4]~22 ));
defparam \result_rb[4]~21 .lut_mask = 16'h96BF;
defparam \result_rb[4]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[5]~23 (
	.dataa(\Add3~7_combout ),
	.datab(\add_in_r_c[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[4]~22 ),
	.combout(\result_rb[5]~23_combout ),
	.cout(\result_rb[5]~24 ));
defparam \result_rb[5]~23 .lut_mask = 16'h96DF;
defparam \result_rb[5]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[6]~25 (
	.dataa(\Add3~6_combout ),
	.datab(\add_in_r_c[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[5]~24 ),
	.combout(\result_rb[6]~25_combout ),
	.cout(\result_rb[6]~26 ));
defparam \result_rb[6]~25 .lut_mask = 16'h96BF;
defparam \result_rb[6]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[7]~27 (
	.dataa(\Add3~5_combout ),
	.datab(\add_in_r_c[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[6]~26 ),
	.combout(\result_rb[7]~27_combout ),
	.cout(\result_rb[7]~28 ));
defparam \result_rb[7]~27 .lut_mask = 16'h96DF;
defparam \result_rb[7]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[8]~29 (
	.dataa(\Add3~4_combout ),
	.datab(\add_in_r_c[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[7]~28 ),
	.combout(\result_rb[8]~29_combout ),
	.cout(\result_rb[8]~30 ));
defparam \result_rb[8]~29 .lut_mask = 16'h96BF;
defparam \result_rb[8]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[9]~31 (
	.dataa(\Add3~3_combout ),
	.datab(\add_in_r_c[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_rb[8]~30 ),
	.combout(\result_rb[9]~31_combout ),
	.cout(\result_rb[9]~32 ));
defparam \result_rb[9]~31 .lut_mask = 16'h96DF;
defparam \result_rb[9]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_rb[10]~33 (
	.dataa(\Add3~3_combout ),
	.datab(\add_in_r_c[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_rb[9]~32 ),
	.combout(\result_rb[10]~33_combout ),
	.cout());
defparam \result_rb[10]~33 .lut_mask = 16'h9696;
defparam \result_rb[10]~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[3]~19 (
	.dataa(\Add1~9_combout ),
	.datab(\add_in_r_a[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[2]~18 ),
	.combout(\result_ra[3]~19_combout ),
	.cout(\result_ra[3]~20 ));
defparam \result_ra[3]~19 .lut_mask = 16'h96DF;
defparam \result_ra[3]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[4]~21 (
	.dataa(\Add1~8_combout ),
	.datab(\add_in_r_a[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[3]~20 ),
	.combout(\result_ra[4]~21_combout ),
	.cout(\result_ra[4]~22 ));
defparam \result_ra[4]~21 .lut_mask = 16'h96BF;
defparam \result_ra[4]~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[5]~23 (
	.dataa(\Add1~7_combout ),
	.datab(\add_in_r_a[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[4]~22 ),
	.combout(\result_ra[5]~23_combout ),
	.cout(\result_ra[5]~24 ));
defparam \result_ra[5]~23 .lut_mask = 16'h96DF;
defparam \result_ra[5]~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[6]~25 (
	.dataa(\Add1~6_combout ),
	.datab(\add_in_r_a[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[5]~24 ),
	.combout(\result_ra[6]~25_combout ),
	.cout(\result_ra[6]~26 ));
defparam \result_ra[6]~25 .lut_mask = 16'h96BF;
defparam \result_ra[6]~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[7]~27 (
	.dataa(\Add1~5_combout ),
	.datab(\add_in_r_a[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[6]~26 ),
	.combout(\result_ra[7]~27_combout ),
	.cout(\result_ra[7]~28 ));
defparam \result_ra[7]~27 .lut_mask = 16'h96DF;
defparam \result_ra[7]~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[8]~29 (
	.dataa(\Add1~4_combout ),
	.datab(\add_in_r_a[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[7]~28 ),
	.combout(\result_ra[8]~29_combout ),
	.cout(\result_ra[8]~30 ));
defparam \result_ra[8]~29 .lut_mask = 16'h96BF;
defparam \result_ra[8]~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[9]~31 (
	.dataa(\Add1~3_combout ),
	.datab(\add_in_r_a[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\result_ra[8]~30 ),
	.combout(\result_ra[9]~31_combout ),
	.cout(\result_ra[9]~32 ));
defparam \result_ra[9]~31 .lut_mask = 16'h96DF;
defparam \result_ra[9]~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \result_ra[10]~33 (
	.dataa(\Add1~3_combout ),
	.datab(\add_in_r_a[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\result_ra[9]~32 ),
	.combout(\result_ra[10]~33_combout ),
	.cout());
defparam \result_ra[10]~33 .lut_mask = 16'h9696;
defparam \result_ra[10]~33 .sum_lutc_input = "cin";

dffeas \offset_counter[8] (
	.clk(clk),
	.d(\offset_counter[8]~26_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[8]~q ),
	.prn(vcc));
defparam \offset_counter[8] .is_wysiwyg = "true";
defparam \offset_counter[8] .power_up = "low";

dffeas \offset_counter[9] (
	.clk(clk),
	.d(\offset_counter[9]~29_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[9]~q ),
	.prn(vcc));
defparam \offset_counter[9] .is_wysiwyg = "true";
defparam \offset_counter[9] .power_up = "low";

dffeas data_val_i(
	.clk(clk),
	.d(\data_val_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\data_val_i~q ),
	.prn(vcc));
defparam data_val_i.is_wysiwyg = "true";
defparam data_val_i.power_up = "low";

dffeas \offset_counter[7] (
	.clk(clk),
	.d(\offset_counter[7]~24_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[7]~q ),
	.prn(vcc));
defparam \offset_counter[7] .is_wysiwyg = "true";
defparam \offset_counter[7] .power_up = "low";

dffeas \offset_counter[6] (
	.clk(clk),
	.d(\offset_counter[6]~22_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[6]~q ),
	.prn(vcc));
defparam \offset_counter[6] .is_wysiwyg = "true";
defparam \offset_counter[6] .power_up = "low";

dffeas \offset_counter[5] (
	.clk(clk),
	.d(\offset_counter[5]~20_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[5]~q ),
	.prn(vcc));
defparam \offset_counter[5] .is_wysiwyg = "true";
defparam \offset_counter[5] .power_up = "low";

dffeas \offset_counter[4] (
	.clk(clk),
	.d(\offset_counter[4]~18_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[4]~q ),
	.prn(vcc));
defparam \offset_counter[4] .is_wysiwyg = "true";
defparam \offset_counter[4] .power_up = "low";

dffeas \offset_counter[3] (
	.clk(clk),
	.d(\offset_counter[3]~16_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[3]~q ),
	.prn(vcc));
defparam \offset_counter[3] .is_wysiwyg = "true";
defparam \offset_counter[3] .power_up = "low";

dffeas \offset_counter[2] (
	.clk(clk),
	.d(\offset_counter[2]~14_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[2]~q ),
	.prn(vcc));
defparam \offset_counter[2] .is_wysiwyg = "true";
defparam \offset_counter[2] .power_up = "low";

dffeas \offset_counter[1] (
	.clk(clk),
	.d(\offset_counter[1]~12_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[1]~q ),
	.prn(vcc));
defparam \offset_counter[1] .is_wysiwyg = "true";
defparam \offset_counter[1] .power_up = "low";

dffeas \offset_counter[0] (
	.clk(clk),
	.d(\offset_counter[0]~10_combout ),
	.asdata(reset_n),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\offset_counter[5]~28_combout ),
	.ena(global_clock_enable),
	.q(\offset_counter[0]~q ),
	.prn(vcc));
defparam \offset_counter[0] .is_wysiwyg = "true";
defparam \offset_counter[0] .power_up = "low";

cycloneive_lcell_comb \offset_counter[0]~10 (
	.dataa(\offset_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\offset_counter[0]~10_combout ),
	.cout(\offset_counter[0]~11 ));
defparam \offset_counter[0]~10 .lut_mask = 16'h55AA;
defparam \offset_counter[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \offset_counter[1]~12 (
	.dataa(\offset_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[0]~11 ),
	.combout(\offset_counter[1]~12_combout ),
	.cout(\offset_counter[1]~13 ));
defparam \offset_counter[1]~12 .lut_mask = 16'h5A5F;
defparam \offset_counter[1]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[2]~14 (
	.dataa(\offset_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[1]~13 ),
	.combout(\offset_counter[2]~14_combout ),
	.cout(\offset_counter[2]~15 ));
defparam \offset_counter[2]~14 .lut_mask = 16'h5AAF;
defparam \offset_counter[2]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[3]~16 (
	.dataa(\offset_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[2]~15 ),
	.combout(\offset_counter[3]~16_combout ),
	.cout(\offset_counter[3]~17 ));
defparam \offset_counter[3]~16 .lut_mask = 16'h5A5F;
defparam \offset_counter[3]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[4]~18 (
	.dataa(\offset_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[3]~17 ),
	.combout(\offset_counter[4]~18_combout ),
	.cout(\offset_counter[4]~19 ));
defparam \offset_counter[4]~18 .lut_mask = 16'h5AAF;
defparam \offset_counter[4]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[5]~20 (
	.dataa(\offset_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[4]~19 ),
	.combout(\offset_counter[5]~20_combout ),
	.cout(\offset_counter[5]~21 ));
defparam \offset_counter[5]~20 .lut_mask = 16'h5A5F;
defparam \offset_counter[5]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[6]~22 (
	.dataa(\offset_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[5]~21 ),
	.combout(\offset_counter[6]~22_combout ),
	.cout(\offset_counter[6]~23 ));
defparam \offset_counter[6]~22 .lut_mask = 16'h5AAF;
defparam \offset_counter[6]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[7]~24 (
	.dataa(\offset_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[6]~23 ),
	.combout(\offset_counter[7]~24_combout ),
	.cout(\offset_counter[7]~25 ));
defparam \offset_counter[7]~24 .lut_mask = 16'h5A5F;
defparam \offset_counter[7]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[8]~26 (
	.dataa(\offset_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\offset_counter[7]~25 ),
	.combout(\offset_counter[8]~26_combout ),
	.cout(\offset_counter[8]~27 ));
defparam \offset_counter[8]~26 .lut_mask = 16'h5AAF;
defparam \offset_counter[8]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \offset_counter[9]~29 (
	.dataa(\offset_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\offset_counter[8]~27 ),
	.combout(\offset_counter[9]~29_combout ),
	.cout());
defparam \offset_counter[9]~29 .lut_mask = 16'h5A5A;
defparam \offset_counter[9]~29 .sum_lutc_input = "cin";

dffeas sgn_2i(
	.clk(clk),
	.d(\sign_vec[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sgn_2i~q ),
	.prn(vcc));
defparam sgn_2i.is_wysiwyg = "true";
defparam sgn_2i.power_up = "low";

cycloneive_lcell_comb \Add11~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[2]~q ),
	.cin(gnd),
	.combout(\Add11~0_combout ),
	.cout());
defparam \Add11~0 .lut_mask = 16'h0FF0;
defparam \Add11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[1]~q ),
	.cin(gnd),
	.combout(\Add11~1_combout ),
	.cout());
defparam \Add11~1 .lut_mask = 16'h0FF0;
defparam \Add11~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[0]~q ),
	.cin(gnd),
	.combout(\Add11~2_combout ),
	.cout());
defparam \Add11~2 .lut_mask = 16'h0FF0;
defparam \Add11~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[10]~q ),
	.cin(gnd),
	.combout(\Add11~3_combout ),
	.cout());
defparam \Add11~3 .lut_mask = 16'h0FF0;
defparam \Add11~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[9]~q ),
	.cin(gnd),
	.combout(\Add11~4_combout ),
	.cout());
defparam \Add11~4 .lut_mask = 16'h0FF0;
defparam \Add11~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[8]~q ),
	.cin(gnd),
	.combout(\Add11~5_combout ),
	.cout());
defparam \Add11~5 .lut_mask = 16'h0FF0;
defparam \Add11~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[7]~q ),
	.cin(gnd),
	.combout(\Add11~6_combout ),
	.cout());
defparam \Add11~6 .lut_mask = 16'h0FF0;
defparam \Add11~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[6]~q ),
	.cin(gnd),
	.combout(\Add11~7_combout ),
	.cout());
defparam \Add11~7 .lut_mask = 16'h0FF0;
defparam \Add11~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[5]~q ),
	.cin(gnd),
	.combout(\Add11~8_combout ),
	.cout());
defparam \Add11~8 .lut_mask = 16'h0FF0;
defparam \Add11~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[4]~q ),
	.cin(gnd),
	.combout(\Add11~9_combout ),
	.cout());
defparam \Add11~9 .lut_mask = 16'h0FF0;
defparam \Add11~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add11~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2i~q ),
	.datad(\result_ib[3]~q ),
	.cin(gnd),
	.combout(\Add11~10_combout ),
	.cout());
defparam \Add11~10 .lut_mask = 16'h0FF0;
defparam \Add11~10 .sum_lutc_input = "datac";

dffeas sgn_2r(
	.clk(clk),
	.d(\sign_vec[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sgn_2r~q ),
	.prn(vcc));
defparam sgn_2r.is_wysiwyg = "true";
defparam sgn_2r.power_up = "low";

cycloneive_lcell_comb \Add9~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[2]~q ),
	.cin(gnd),
	.combout(\Add9~0_combout ),
	.cout());
defparam \Add9~0 .lut_mask = 16'h0FF0;
defparam \Add9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[1]~q ),
	.cin(gnd),
	.combout(\Add9~1_combout ),
	.cout());
defparam \Add9~1 .lut_mask = 16'h0FF0;
defparam \Add9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[0]~q ),
	.cin(gnd),
	.combout(\Add9~2_combout ),
	.cout());
defparam \Add9~2 .lut_mask = 16'h0FF0;
defparam \Add9~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[10]~q ),
	.cin(gnd),
	.combout(\Add9~3_combout ),
	.cout());
defparam \Add9~3 .lut_mask = 16'h0FF0;
defparam \Add9~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[9]~q ),
	.cin(gnd),
	.combout(\Add9~4_combout ),
	.cout());
defparam \Add9~4 .lut_mask = 16'h0FF0;
defparam \Add9~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[8]~q ),
	.cin(gnd),
	.combout(\Add9~5_combout ),
	.cout());
defparam \Add9~5 .lut_mask = 16'h0FF0;
defparam \Add9~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[7]~q ),
	.cin(gnd),
	.combout(\Add9~6_combout ),
	.cout());
defparam \Add9~6 .lut_mask = 16'h0FF0;
defparam \Add9~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[6]~q ),
	.cin(gnd),
	.combout(\Add9~7_combout ),
	.cout());
defparam \Add9~7 .lut_mask = 16'h0FF0;
defparam \Add9~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[5]~q ),
	.cin(gnd),
	.combout(\Add9~8_combout ),
	.cout());
defparam \Add9~8 .lut_mask = 16'h0FF0;
defparam \Add9~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[4]~q ),
	.cin(gnd),
	.combout(\Add9~9_combout ),
	.cout());
defparam \Add9~9 .lut_mask = 16'h0FF0;
defparam \Add9~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add9~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sgn_2r~q ),
	.datad(\result_rb[3]~q ),
	.cin(gnd),
	.combout(\Add9~10_combout ),
	.cout());
defparam \Add9~10 .lut_mask = 16'h0FF0;
defparam \Add9~10 .sum_lutc_input = "datac";

dffeas \sign_vec[0] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_vec[0]~q ),
	.prn(vcc));
defparam \sign_vec[0] .is_wysiwyg = "true";
defparam \sign_vec[0] .power_up = "low";

dffeas \add_in_i_d[2] (
	.clk(clk),
	.d(\add_in_i_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[2]~q ),
	.prn(vcc));
defparam \add_in_i_d[2] .is_wysiwyg = "true";
defparam \add_in_i_d[2] .power_up = "low";

dffeas \sign_vec[3] (
	.clk(clk),
	.d(\sign_vec[3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_vec[3]~q ),
	.prn(vcc));
defparam \sign_vec[3] .is_wysiwyg = "true";
defparam \sign_vec[3] .power_up = "low";

cycloneive_lcell_comb \Add4~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\add_in_i_d[2]~q ),
	.datad(\sign_vec[3]~q ),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout());
defparam \Add4~0 .lut_mask = 16'h0FF0;
defparam \Add4~0 .sum_lutc_input = "datac";

dffeas \add_in_i_c[2] (
	.clk(clk),
	.d(\add_in_i_c~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[2]~q ),
	.prn(vcc));
defparam \add_in_i_c[2] .is_wysiwyg = "true";
defparam \add_in_i_c[2] .power_up = "low";

dffeas \add_in_i_d[1] (
	.clk(clk),
	.d(\add_in_i_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[1]~q ),
	.prn(vcc));
defparam \add_in_i_d[1] .is_wysiwyg = "true";
defparam \add_in_i_d[1] .power_up = "low";

cycloneive_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[1]~q ),
	.cin(gnd),
	.combout(\Add4~1_combout ),
	.cout());
defparam \Add4~1 .lut_mask = 16'h0FF0;
defparam \Add4~1 .sum_lutc_input = "datac";

dffeas \add_in_i_c[1] (
	.clk(clk),
	.d(\add_in_i_c~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[1]~q ),
	.prn(vcc));
defparam \add_in_i_c[1] .is_wysiwyg = "true";
defparam \add_in_i_c[1] .power_up = "low";

dffeas \add_in_i_d[0] (
	.clk(clk),
	.d(\add_in_i_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[0]~q ),
	.prn(vcc));
defparam \add_in_i_d[0] .is_wysiwyg = "true";
defparam \add_in_i_d[0] .power_up = "low";

cycloneive_lcell_comb \Add4~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[0]~q ),
	.cin(gnd),
	.combout(\Add4~2_combout ),
	.cout());
defparam \Add4~2 .lut_mask = 16'h0FF0;
defparam \Add4~2 .sum_lutc_input = "datac";

dffeas \add_in_i_c[0] (
	.clk(clk),
	.d(\add_in_i_c~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[0]~q ),
	.prn(vcc));
defparam \add_in_i_c[0] .is_wysiwyg = "true";
defparam \add_in_i_c[0] .power_up = "low";

dffeas \add_in_i_b[2] (
	.clk(clk),
	.d(data_3_imag_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[2]~q ),
	.prn(vcc));
defparam \add_in_i_b[2] .is_wysiwyg = "true";
defparam \add_in_i_b[2] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[2]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h0FF0;
defparam \Add2~0 .sum_lutc_input = "datac";

dffeas \add_in_i_a[2] (
	.clk(clk),
	.d(data_1_imag_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[2]~q ),
	.prn(vcc));
defparam \add_in_i_a[2] .is_wysiwyg = "true";
defparam \add_in_i_a[2] .power_up = "low";

dffeas \add_in_i_b[1] (
	.clk(clk),
	.d(data_3_imag_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[1]~q ),
	.prn(vcc));
defparam \add_in_i_b[1] .is_wysiwyg = "true";
defparam \add_in_i_b[1] .power_up = "low";

cycloneive_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[1]~q ),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h0FF0;
defparam \Add2~1 .sum_lutc_input = "datac";

dffeas \add_in_i_a[1] (
	.clk(clk),
	.d(data_1_imag_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[1]~q ),
	.prn(vcc));
defparam \add_in_i_a[1] .is_wysiwyg = "true";
defparam \add_in_i_a[1] .power_up = "low";

dffeas \add_in_i_b[0] (
	.clk(clk),
	.d(data_3_imag_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[0]~q ),
	.prn(vcc));
defparam \add_in_i_b[0] .is_wysiwyg = "true";
defparam \add_in_i_b[0] .power_up = "low";

cycloneive_lcell_comb \Add2~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[0]~q ),
	.cin(gnd),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h0FF0;
defparam \Add2~2 .sum_lutc_input = "datac";

dffeas \add_in_i_a[0] (
	.clk(clk),
	.d(data_1_imag_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[0]~q ),
	.prn(vcc));
defparam \add_in_i_a[0] .is_wysiwyg = "true";
defparam \add_in_i_a[0] .power_up = "low";

dffeas \add_in_i_d[9] (
	.clk(clk),
	.d(\add_in_i_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[9]~q ),
	.prn(vcc));
defparam \add_in_i_d[9] .is_wysiwyg = "true";
defparam \add_in_i_d[9] .power_up = "low";

cycloneive_lcell_comb \Add4~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[9]~q ),
	.cin(gnd),
	.combout(\Add4~3_combout ),
	.cout());
defparam \Add4~3 .lut_mask = 16'h0FF0;
defparam \Add4~3 .sum_lutc_input = "datac";

dffeas \add_in_i_c[9] (
	.clk(clk),
	.d(\add_in_i_c~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[9]~q ),
	.prn(vcc));
defparam \add_in_i_c[9] .is_wysiwyg = "true";
defparam \add_in_i_c[9] .power_up = "low";

dffeas \add_in_i_d[8] (
	.clk(clk),
	.d(\add_in_i_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[8]~q ),
	.prn(vcc));
defparam \add_in_i_d[8] .is_wysiwyg = "true";
defparam \add_in_i_d[8] .power_up = "low";

cycloneive_lcell_comb \Add4~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[8]~q ),
	.cin(gnd),
	.combout(\Add4~4_combout ),
	.cout());
defparam \Add4~4 .lut_mask = 16'h0FF0;
defparam \Add4~4 .sum_lutc_input = "datac";

dffeas \add_in_i_c[8] (
	.clk(clk),
	.d(\add_in_i_c~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[8]~q ),
	.prn(vcc));
defparam \add_in_i_c[8] .is_wysiwyg = "true";
defparam \add_in_i_c[8] .power_up = "low";

dffeas \add_in_i_d[7] (
	.clk(clk),
	.d(\add_in_i_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[7]~q ),
	.prn(vcc));
defparam \add_in_i_d[7] .is_wysiwyg = "true";
defparam \add_in_i_d[7] .power_up = "low";

cycloneive_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[7]~q ),
	.cin(gnd),
	.combout(\Add4~5_combout ),
	.cout());
defparam \Add4~5 .lut_mask = 16'h0FF0;
defparam \Add4~5 .sum_lutc_input = "datac";

dffeas \add_in_i_c[7] (
	.clk(clk),
	.d(\add_in_i_c~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[7]~q ),
	.prn(vcc));
defparam \add_in_i_c[7] .is_wysiwyg = "true";
defparam \add_in_i_c[7] .power_up = "low";

dffeas \add_in_i_d[6] (
	.clk(clk),
	.d(\add_in_i_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[6]~q ),
	.prn(vcc));
defparam \add_in_i_d[6] .is_wysiwyg = "true";
defparam \add_in_i_d[6] .power_up = "low";

cycloneive_lcell_comb \Add4~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[6]~q ),
	.cin(gnd),
	.combout(\Add4~6_combout ),
	.cout());
defparam \Add4~6 .lut_mask = 16'h0FF0;
defparam \Add4~6 .sum_lutc_input = "datac";

dffeas \add_in_i_c[6] (
	.clk(clk),
	.d(\add_in_i_c~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[6]~q ),
	.prn(vcc));
defparam \add_in_i_c[6] .is_wysiwyg = "true";
defparam \add_in_i_c[6] .power_up = "low";

dffeas \add_in_i_d[5] (
	.clk(clk),
	.d(\add_in_i_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[5]~q ),
	.prn(vcc));
defparam \add_in_i_d[5] .is_wysiwyg = "true";
defparam \add_in_i_d[5] .power_up = "low";

cycloneive_lcell_comb \Add4~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[5]~q ),
	.cin(gnd),
	.combout(\Add4~7_combout ),
	.cout());
defparam \Add4~7 .lut_mask = 16'h0FF0;
defparam \Add4~7 .sum_lutc_input = "datac";

dffeas \add_in_i_c[5] (
	.clk(clk),
	.d(\add_in_i_c~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[5]~q ),
	.prn(vcc));
defparam \add_in_i_c[5] .is_wysiwyg = "true";
defparam \add_in_i_c[5] .power_up = "low";

dffeas \add_in_i_d[4] (
	.clk(clk),
	.d(\add_in_i_d~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[4]~q ),
	.prn(vcc));
defparam \add_in_i_d[4] .is_wysiwyg = "true";
defparam \add_in_i_d[4] .power_up = "low";

cycloneive_lcell_comb \Add4~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[4]~q ),
	.cin(gnd),
	.combout(\Add4~8_combout ),
	.cout());
defparam \Add4~8 .lut_mask = 16'h0FF0;
defparam \Add4~8 .sum_lutc_input = "datac";

dffeas \add_in_i_c[4] (
	.clk(clk),
	.d(\add_in_i_c~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[4]~q ),
	.prn(vcc));
defparam \add_in_i_c[4] .is_wysiwyg = "true";
defparam \add_in_i_c[4] .power_up = "low";

dffeas \add_in_i_d[3] (
	.clk(clk),
	.d(\add_in_i_d~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_d[3]~q ),
	.prn(vcc));
defparam \add_in_i_d[3] .is_wysiwyg = "true";
defparam \add_in_i_d[3] .power_up = "low";

cycloneive_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_d[3]~q ),
	.cin(gnd),
	.combout(\Add4~9_combout ),
	.cout());
defparam \Add4~9 .lut_mask = 16'h0FF0;
defparam \Add4~9 .sum_lutc_input = "datac";

dffeas \add_in_i_c[3] (
	.clk(clk),
	.d(\add_in_i_c~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_c[3]~q ),
	.prn(vcc));
defparam \add_in_i_c[3] .is_wysiwyg = "true";
defparam \add_in_i_c[3] .power_up = "low";

dffeas \add_in_i_b[9] (
	.clk(clk),
	.d(data_3_imag_i[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[9]~q ),
	.prn(vcc));
defparam \add_in_i_b[9] .is_wysiwyg = "true";
defparam \add_in_i_b[9] .power_up = "low";

cycloneive_lcell_comb \Add2~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[9]~q ),
	.cin(gnd),
	.combout(\Add2~3_combout ),
	.cout());
defparam \Add2~3 .lut_mask = 16'h0FF0;
defparam \Add2~3 .sum_lutc_input = "datac";

dffeas \add_in_i_a[9] (
	.clk(clk),
	.d(data_1_imag_i[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[9]~q ),
	.prn(vcc));
defparam \add_in_i_a[9] .is_wysiwyg = "true";
defparam \add_in_i_a[9] .power_up = "low";

dffeas \add_in_i_b[8] (
	.clk(clk),
	.d(data_3_imag_i[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[8]~q ),
	.prn(vcc));
defparam \add_in_i_b[8] .is_wysiwyg = "true";
defparam \add_in_i_b[8] .power_up = "low";

cycloneive_lcell_comb \Add2~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[8]~q ),
	.cin(gnd),
	.combout(\Add2~4_combout ),
	.cout());
defparam \Add2~4 .lut_mask = 16'h0FF0;
defparam \Add2~4 .sum_lutc_input = "datac";

dffeas \add_in_i_a[8] (
	.clk(clk),
	.d(data_1_imag_i[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[8]~q ),
	.prn(vcc));
defparam \add_in_i_a[8] .is_wysiwyg = "true";
defparam \add_in_i_a[8] .power_up = "low";

dffeas \add_in_i_b[7] (
	.clk(clk),
	.d(data_3_imag_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[7]~q ),
	.prn(vcc));
defparam \add_in_i_b[7] .is_wysiwyg = "true";
defparam \add_in_i_b[7] .power_up = "low";

cycloneive_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[7]~q ),
	.cin(gnd),
	.combout(\Add2~5_combout ),
	.cout());
defparam \Add2~5 .lut_mask = 16'h0FF0;
defparam \Add2~5 .sum_lutc_input = "datac";

dffeas \add_in_i_a[7] (
	.clk(clk),
	.d(data_1_imag_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[7]~q ),
	.prn(vcc));
defparam \add_in_i_a[7] .is_wysiwyg = "true";
defparam \add_in_i_a[7] .power_up = "low";

dffeas \add_in_i_b[6] (
	.clk(clk),
	.d(data_3_imag_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[6]~q ),
	.prn(vcc));
defparam \add_in_i_b[6] .is_wysiwyg = "true";
defparam \add_in_i_b[6] .power_up = "low";

cycloneive_lcell_comb \Add2~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[6]~q ),
	.cin(gnd),
	.combout(\Add2~6_combout ),
	.cout());
defparam \Add2~6 .lut_mask = 16'h0FF0;
defparam \Add2~6 .sum_lutc_input = "datac";

dffeas \add_in_i_a[6] (
	.clk(clk),
	.d(data_1_imag_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[6]~q ),
	.prn(vcc));
defparam \add_in_i_a[6] .is_wysiwyg = "true";
defparam \add_in_i_a[6] .power_up = "low";

dffeas \add_in_i_b[5] (
	.clk(clk),
	.d(data_3_imag_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[5]~q ),
	.prn(vcc));
defparam \add_in_i_b[5] .is_wysiwyg = "true";
defparam \add_in_i_b[5] .power_up = "low";

cycloneive_lcell_comb \Add2~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[5]~q ),
	.cin(gnd),
	.combout(\Add2~7_combout ),
	.cout());
defparam \Add2~7 .lut_mask = 16'h0FF0;
defparam \Add2~7 .sum_lutc_input = "datac";

dffeas \add_in_i_a[5] (
	.clk(clk),
	.d(data_1_imag_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[5]~q ),
	.prn(vcc));
defparam \add_in_i_a[5] .is_wysiwyg = "true";
defparam \add_in_i_a[5] .power_up = "low";

dffeas \add_in_i_b[4] (
	.clk(clk),
	.d(data_3_imag_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[4]~q ),
	.prn(vcc));
defparam \add_in_i_b[4] .is_wysiwyg = "true";
defparam \add_in_i_b[4] .power_up = "low";

cycloneive_lcell_comb \Add2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[4]~q ),
	.cin(gnd),
	.combout(\Add2~8_combout ),
	.cout());
defparam \Add2~8 .lut_mask = 16'h0FF0;
defparam \Add2~8 .sum_lutc_input = "datac";

dffeas \add_in_i_a[4] (
	.clk(clk),
	.d(data_1_imag_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[4]~q ),
	.prn(vcc));
defparam \add_in_i_a[4] .is_wysiwyg = "true";
defparam \add_in_i_a[4] .power_up = "low";

dffeas \add_in_i_b[3] (
	.clk(clk),
	.d(data_3_imag_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_b[3]~q ),
	.prn(vcc));
defparam \add_in_i_b[3] .is_wysiwyg = "true";
defparam \add_in_i_b[3] .power_up = "low";

cycloneive_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_i_b[3]~q ),
	.cin(gnd),
	.combout(\Add2~9_combout ),
	.cout());
defparam \Add2~9 .lut_mask = 16'h0FF0;
defparam \Add2~9 .sum_lutc_input = "datac";

dffeas \add_in_i_a[3] (
	.clk(clk),
	.d(data_1_imag_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_i_a[3]~q ),
	.prn(vcc));
defparam \add_in_i_a[3] .is_wysiwyg = "true";
defparam \add_in_i_a[3] .power_up = "low";

dffeas \sign_vec[1] (
	.clk(clk),
	.d(\sign_vec[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_vec[1]~q ),
	.prn(vcc));
defparam \sign_vec[1] .is_wysiwyg = "true";
defparam \sign_vec[1] .power_up = "low";

dffeas \add_in_r_d[2] (
	.clk(clk),
	.d(\add_in_r_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[2]~q ),
	.prn(vcc));
defparam \add_in_r_d[2] .is_wysiwyg = "true";
defparam \add_in_r_d[2] .power_up = "low";

cycloneive_lcell_comb \Add3~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[2]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h0FF0;
defparam \Add3~0 .sum_lutc_input = "datac";

dffeas \add_in_r_c[2] (
	.clk(clk),
	.d(\add_in_r_c~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[2]~q ),
	.prn(vcc));
defparam \add_in_r_c[2] .is_wysiwyg = "true";
defparam \add_in_r_c[2] .power_up = "low";

dffeas \add_in_r_d[1] (
	.clk(clk),
	.d(\add_in_r_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[1]~q ),
	.prn(vcc));
defparam \add_in_r_d[1] .is_wysiwyg = "true";
defparam \add_in_r_d[1] .power_up = "low";

cycloneive_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[1]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'h0FF0;
defparam \Add3~1 .sum_lutc_input = "datac";

dffeas \add_in_r_c[1] (
	.clk(clk),
	.d(\add_in_r_c~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[1]~q ),
	.prn(vcc));
defparam \add_in_r_c[1] .is_wysiwyg = "true";
defparam \add_in_r_c[1] .power_up = "low";

dffeas \add_in_r_d[0] (
	.clk(clk),
	.d(\add_in_r_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[0]~q ),
	.prn(vcc));
defparam \add_in_r_d[0] .is_wysiwyg = "true";
defparam \add_in_r_d[0] .power_up = "low";

cycloneive_lcell_comb \Add3~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[0]~q ),
	.cin(gnd),
	.combout(\Add3~2_combout ),
	.cout());
defparam \Add3~2 .lut_mask = 16'h0FF0;
defparam \Add3~2 .sum_lutc_input = "datac";

dffeas \add_in_r_c[0] (
	.clk(clk),
	.d(\add_in_r_c~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[0]~q ),
	.prn(vcc));
defparam \add_in_r_c[0] .is_wysiwyg = "true";
defparam \add_in_r_c[0] .power_up = "low";

dffeas \add_in_r_b[2] (
	.clk(clk),
	.d(data_3_real_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[2]~q ),
	.prn(vcc));
defparam \add_in_r_b[2] .is_wysiwyg = "true";
defparam \add_in_r_b[2] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[2]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas \add_in_r_a[2] (
	.clk(clk),
	.d(data_1_real_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[2]~q ),
	.prn(vcc));
defparam \add_in_r_a[2] .is_wysiwyg = "true";
defparam \add_in_r_a[2] .power_up = "low";

dffeas \add_in_r_b[1] (
	.clk(clk),
	.d(data_3_real_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[1]~q ),
	.prn(vcc));
defparam \add_in_r_b[1] .is_wysiwyg = "true";
defparam \add_in_r_b[1] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[1]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

dffeas \add_in_r_a[1] (
	.clk(clk),
	.d(data_1_real_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[1]~q ),
	.prn(vcc));
defparam \add_in_r_a[1] .is_wysiwyg = "true";
defparam \add_in_r_a[1] .power_up = "low";

dffeas \add_in_r_b[0] (
	.clk(clk),
	.d(data_3_real_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[0]~q ),
	.prn(vcc));
defparam \add_in_r_b[0] .is_wysiwyg = "true";
defparam \add_in_r_b[0] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[0]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

dffeas \add_in_r_a[0] (
	.clk(clk),
	.d(data_1_real_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[0]~q ),
	.prn(vcc));
defparam \add_in_r_a[0] .is_wysiwyg = "true";
defparam \add_in_r_a[0] .power_up = "low";

dffeas \add_in_r_d[9] (
	.clk(clk),
	.d(\add_in_r_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[9]~q ),
	.prn(vcc));
defparam \add_in_r_d[9] .is_wysiwyg = "true";
defparam \add_in_r_d[9] .power_up = "low";

cycloneive_lcell_comb \Add3~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[9]~q ),
	.cin(gnd),
	.combout(\Add3~3_combout ),
	.cout());
defparam \Add3~3 .lut_mask = 16'h0FF0;
defparam \Add3~3 .sum_lutc_input = "datac";

dffeas \add_in_r_c[9] (
	.clk(clk),
	.d(\add_in_r_c~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[9]~q ),
	.prn(vcc));
defparam \add_in_r_c[9] .is_wysiwyg = "true";
defparam \add_in_r_c[9] .power_up = "low";

dffeas \add_in_r_d[8] (
	.clk(clk),
	.d(\add_in_r_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[8]~q ),
	.prn(vcc));
defparam \add_in_r_d[8] .is_wysiwyg = "true";
defparam \add_in_r_d[8] .power_up = "low";

cycloneive_lcell_comb \Add3~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[8]~q ),
	.cin(gnd),
	.combout(\Add3~4_combout ),
	.cout());
defparam \Add3~4 .lut_mask = 16'h0FF0;
defparam \Add3~4 .sum_lutc_input = "datac";

dffeas \add_in_r_c[8] (
	.clk(clk),
	.d(\add_in_r_c~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[8]~q ),
	.prn(vcc));
defparam \add_in_r_c[8] .is_wysiwyg = "true";
defparam \add_in_r_c[8] .power_up = "low";

dffeas \add_in_r_d[7] (
	.clk(clk),
	.d(\add_in_r_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[7]~q ),
	.prn(vcc));
defparam \add_in_r_d[7] .is_wysiwyg = "true";
defparam \add_in_r_d[7] .power_up = "low";

cycloneive_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[7]~q ),
	.cin(gnd),
	.combout(\Add3~5_combout ),
	.cout());
defparam \Add3~5 .lut_mask = 16'h0FF0;
defparam \Add3~5 .sum_lutc_input = "datac";

dffeas \add_in_r_c[7] (
	.clk(clk),
	.d(\add_in_r_c~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[7]~q ),
	.prn(vcc));
defparam \add_in_r_c[7] .is_wysiwyg = "true";
defparam \add_in_r_c[7] .power_up = "low";

dffeas \add_in_r_d[6] (
	.clk(clk),
	.d(\add_in_r_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[6]~q ),
	.prn(vcc));
defparam \add_in_r_d[6] .is_wysiwyg = "true";
defparam \add_in_r_d[6] .power_up = "low";

cycloneive_lcell_comb \Add3~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[6]~q ),
	.cin(gnd),
	.combout(\Add3~6_combout ),
	.cout());
defparam \Add3~6 .lut_mask = 16'h0FF0;
defparam \Add3~6 .sum_lutc_input = "datac";

dffeas \add_in_r_c[6] (
	.clk(clk),
	.d(\add_in_r_c~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[6]~q ),
	.prn(vcc));
defparam \add_in_r_c[6] .is_wysiwyg = "true";
defparam \add_in_r_c[6] .power_up = "low";

dffeas \add_in_r_d[5] (
	.clk(clk),
	.d(\add_in_r_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[5]~q ),
	.prn(vcc));
defparam \add_in_r_d[5] .is_wysiwyg = "true";
defparam \add_in_r_d[5] .power_up = "low";

cycloneive_lcell_comb \Add3~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[5]~q ),
	.cin(gnd),
	.combout(\Add3~7_combout ),
	.cout());
defparam \Add3~7 .lut_mask = 16'h0FF0;
defparam \Add3~7 .sum_lutc_input = "datac";

dffeas \add_in_r_c[5] (
	.clk(clk),
	.d(\add_in_r_c~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[5]~q ),
	.prn(vcc));
defparam \add_in_r_c[5] .is_wysiwyg = "true";
defparam \add_in_r_c[5] .power_up = "low";

dffeas \add_in_r_d[4] (
	.clk(clk),
	.d(\add_in_r_d~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[4]~q ),
	.prn(vcc));
defparam \add_in_r_d[4] .is_wysiwyg = "true";
defparam \add_in_r_d[4] .power_up = "low";

cycloneive_lcell_comb \Add3~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[4]~q ),
	.cin(gnd),
	.combout(\Add3~8_combout ),
	.cout());
defparam \Add3~8 .lut_mask = 16'h0FF0;
defparam \Add3~8 .sum_lutc_input = "datac";

dffeas \add_in_r_c[4] (
	.clk(clk),
	.d(\add_in_r_c~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[4]~q ),
	.prn(vcc));
defparam \add_in_r_c[4] .is_wysiwyg = "true";
defparam \add_in_r_c[4] .power_up = "low";

dffeas \add_in_r_d[3] (
	.clk(clk),
	.d(\add_in_r_d~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_d[3]~q ),
	.prn(vcc));
defparam \add_in_r_d[3] .is_wysiwyg = "true";
defparam \add_in_r_d[3] .power_up = "low";

cycloneive_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_d[3]~q ),
	.cin(gnd),
	.combout(\Add3~9_combout ),
	.cout());
defparam \Add3~9 .lut_mask = 16'h0FF0;
defparam \Add3~9 .sum_lutc_input = "datac";

dffeas \add_in_r_c[3] (
	.clk(clk),
	.d(\add_in_r_c~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_c[3]~q ),
	.prn(vcc));
defparam \add_in_r_c[3] .is_wysiwyg = "true";
defparam \add_in_r_c[3] .power_up = "low";

dffeas \add_in_r_b[9] (
	.clk(clk),
	.d(data_3_real_i[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[9]~q ),
	.prn(vcc));
defparam \add_in_r_b[9] .is_wysiwyg = "true";
defparam \add_in_r_b[9] .power_up = "low";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[9]~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

dffeas \add_in_r_a[9] (
	.clk(clk),
	.d(data_1_real_i[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[9]~q ),
	.prn(vcc));
defparam \add_in_r_a[9] .is_wysiwyg = "true";
defparam \add_in_r_a[9] .power_up = "low";

dffeas \add_in_r_b[8] (
	.clk(clk),
	.d(data_3_real_i[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[8]~q ),
	.prn(vcc));
defparam \add_in_r_b[8] .is_wysiwyg = "true";
defparam \add_in_r_b[8] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[8]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

dffeas \add_in_r_a[8] (
	.clk(clk),
	.d(data_1_real_i[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[8]~q ),
	.prn(vcc));
defparam \add_in_r_a[8] .is_wysiwyg = "true";
defparam \add_in_r_a[8] .power_up = "low";

dffeas \add_in_r_b[7] (
	.clk(clk),
	.d(data_3_real_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[7]~q ),
	.prn(vcc));
defparam \add_in_r_b[7] .is_wysiwyg = "true";
defparam \add_in_r_b[7] .power_up = "low";

cycloneive_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[7]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

dffeas \add_in_r_a[7] (
	.clk(clk),
	.d(data_1_real_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[7]~q ),
	.prn(vcc));
defparam \add_in_r_a[7] .is_wysiwyg = "true";
defparam \add_in_r_a[7] .power_up = "low";

dffeas \add_in_r_b[6] (
	.clk(clk),
	.d(data_3_real_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[6]~q ),
	.prn(vcc));
defparam \add_in_r_b[6] .is_wysiwyg = "true";
defparam \add_in_r_b[6] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[6]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

dffeas \add_in_r_a[6] (
	.clk(clk),
	.d(data_1_real_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[6]~q ),
	.prn(vcc));
defparam \add_in_r_a[6] .is_wysiwyg = "true";
defparam \add_in_r_a[6] .power_up = "low";

dffeas \add_in_r_b[5] (
	.clk(clk),
	.d(data_3_real_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[5]~q ),
	.prn(vcc));
defparam \add_in_r_b[5] .is_wysiwyg = "true";
defparam \add_in_r_b[5] .power_up = "low";

cycloneive_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[5]~q ),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

dffeas \add_in_r_a[5] (
	.clk(clk),
	.d(data_1_real_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[5]~q ),
	.prn(vcc));
defparam \add_in_r_a[5] .is_wysiwyg = "true";
defparam \add_in_r_a[5] .power_up = "low";

dffeas \add_in_r_b[4] (
	.clk(clk),
	.d(data_3_real_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[4]~q ),
	.prn(vcc));
defparam \add_in_r_b[4] .is_wysiwyg = "true";
defparam \add_in_r_b[4] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[4]~q ),
	.cin(gnd),
	.combout(\Add1~8_combout ),
	.cout());
defparam \Add1~8 .lut_mask = 16'h0FF0;
defparam \Add1~8 .sum_lutc_input = "datac";

dffeas \add_in_r_a[4] (
	.clk(clk),
	.d(data_1_real_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[4]~q ),
	.prn(vcc));
defparam \add_in_r_a[4] .is_wysiwyg = "true";
defparam \add_in_r_a[4] .power_up = "low";

dffeas \add_in_r_b[3] (
	.clk(clk),
	.d(data_3_real_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_b[3]~q ),
	.prn(vcc));
defparam \add_in_r_b[3] .is_wysiwyg = "true";
defparam \add_in_r_b[3] .power_up = "low";

cycloneive_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_vec[3]~q ),
	.datad(\add_in_r_b[3]~q ),
	.cin(gnd),
	.combout(\Add1~9_combout ),
	.cout());
defparam \Add1~9 .lut_mask = 16'h0FF0;
defparam \Add1~9 .sum_lutc_input = "datac";

dffeas \add_in_r_a[3] (
	.clk(clk),
	.d(data_1_real_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\add_in_r_a[3]~q ),
	.prn(vcc));
defparam \add_in_r_a[3] .is_wysiwyg = "true";
defparam \add_in_r_a[3] .power_up = "low";

dffeas \sign_sel[0] (
	.clk(clk),
	.d(\offset_counter[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_sel[0]~q ),
	.prn(vcc));
defparam \sign_sel[0] .is_wysiwyg = "true";
defparam \sign_sel[0] .power_up = "low";

dffeas \sign_sel[1] (
	.clk(clk),
	.d(\offset_counter[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\sign_sel[1]~q ),
	.prn(vcc));
defparam \sign_sel[1] .is_wysiwyg = "true";
defparam \sign_sel[1] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sign_sel[0]~q ),
	.datad(\sign_sel[1]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h0FF0;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~0 (
	.dataa(ram_in_reg_2_3),
	.datab(ram_in_reg_2_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~0_combout ),
	.cout());
defparam \add_in_i_d~0 .lut_mask = 16'hAACC;
defparam \add_in_i_d~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~0 (
	.dataa(ram_in_reg_2_1),
	.datab(ram_in_reg_2_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~0_combout ),
	.cout());
defparam \add_in_i_c~0 .lut_mask = 16'hAACC;
defparam \add_in_i_c~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~1 (
	.dataa(ram_in_reg_1_3),
	.datab(ram_in_reg_1_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~1_combout ),
	.cout());
defparam \add_in_i_d~1 .lut_mask = 16'hAACC;
defparam \add_in_i_d~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~1 (
	.dataa(ram_in_reg_1_1),
	.datab(ram_in_reg_1_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~1_combout ),
	.cout());
defparam \add_in_i_c~1 .lut_mask = 16'hAACC;
defparam \add_in_i_c~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~2 (
	.dataa(ram_in_reg_0_3),
	.datab(ram_in_reg_0_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~2_combout ),
	.cout());
defparam \add_in_i_d~2 .lut_mask = 16'hAACC;
defparam \add_in_i_d~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~2 (
	.dataa(ram_in_reg_0_1),
	.datab(ram_in_reg_0_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~2_combout ),
	.cout());
defparam \add_in_i_c~2 .lut_mask = 16'hAACC;
defparam \add_in_i_c~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~3 (
	.dataa(ram_in_reg_9_3),
	.datab(ram_in_reg_9_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~3_combout ),
	.cout());
defparam \add_in_i_d~3 .lut_mask = 16'hAACC;
defparam \add_in_i_d~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~3 (
	.dataa(ram_in_reg_9_1),
	.datab(ram_in_reg_9_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~3_combout ),
	.cout());
defparam \add_in_i_c~3 .lut_mask = 16'hAACC;
defparam \add_in_i_c~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~4 (
	.dataa(ram_in_reg_8_3),
	.datab(ram_in_reg_8_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~4_combout ),
	.cout());
defparam \add_in_i_d~4 .lut_mask = 16'hAACC;
defparam \add_in_i_d~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~4 (
	.dataa(ram_in_reg_8_1),
	.datab(ram_in_reg_8_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~4_combout ),
	.cout());
defparam \add_in_i_c~4 .lut_mask = 16'hAACC;
defparam \add_in_i_c~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~5 (
	.dataa(ram_in_reg_7_3),
	.datab(ram_in_reg_7_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~5_combout ),
	.cout());
defparam \add_in_i_d~5 .lut_mask = 16'hAACC;
defparam \add_in_i_d~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~5 (
	.dataa(ram_in_reg_7_1),
	.datab(ram_in_reg_7_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~5_combout ),
	.cout());
defparam \add_in_i_c~5 .lut_mask = 16'hAACC;
defparam \add_in_i_c~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~6 (
	.dataa(ram_in_reg_6_3),
	.datab(ram_in_reg_6_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~6_combout ),
	.cout());
defparam \add_in_i_d~6 .lut_mask = 16'hAACC;
defparam \add_in_i_d~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~6 (
	.dataa(ram_in_reg_6_1),
	.datab(ram_in_reg_6_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~6_combout ),
	.cout());
defparam \add_in_i_c~6 .lut_mask = 16'hAACC;
defparam \add_in_i_c~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~7 (
	.dataa(ram_in_reg_5_3),
	.datab(ram_in_reg_5_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~7_combout ),
	.cout());
defparam \add_in_i_d~7 .lut_mask = 16'hAACC;
defparam \add_in_i_d~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~7 (
	.dataa(ram_in_reg_5_1),
	.datab(ram_in_reg_5_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~7_combout ),
	.cout());
defparam \add_in_i_c~7 .lut_mask = 16'hAACC;
defparam \add_in_i_c~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~8 (
	.dataa(ram_in_reg_4_3),
	.datab(ram_in_reg_4_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~8_combout ),
	.cout());
defparam \add_in_i_d~8 .lut_mask = 16'hAACC;
defparam \add_in_i_d~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~8 (
	.dataa(ram_in_reg_4_1),
	.datab(ram_in_reg_4_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~8_combout ),
	.cout());
defparam \add_in_i_c~8 .lut_mask = 16'hAACC;
defparam \add_in_i_c~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_d~9 (
	.dataa(ram_in_reg_3_3),
	.datab(ram_in_reg_3_7),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_d~9_combout ),
	.cout());
defparam \add_in_i_d~9 .lut_mask = 16'hAACC;
defparam \add_in_i_d~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_i_c~9 (
	.dataa(ram_in_reg_3_1),
	.datab(ram_in_reg_3_5),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_i_c~9_combout ),
	.cout());
defparam \add_in_i_c~9 .lut_mask = 16'hAACC;
defparam \add_in_i_c~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~0 (
	.dataa(ram_in_reg_2_7),
	.datab(ram_in_reg_2_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~0_combout ),
	.cout());
defparam \add_in_r_d~0 .lut_mask = 16'hAACC;
defparam \add_in_r_d~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~0 (
	.dataa(ram_in_reg_2_5),
	.datab(ram_in_reg_2_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~0_combout ),
	.cout());
defparam \add_in_r_c~0 .lut_mask = 16'hAACC;
defparam \add_in_r_c~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~1 (
	.dataa(ram_in_reg_1_7),
	.datab(ram_in_reg_1_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~1_combout ),
	.cout());
defparam \add_in_r_d~1 .lut_mask = 16'hAACC;
defparam \add_in_r_d~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~1 (
	.dataa(ram_in_reg_1_5),
	.datab(ram_in_reg_1_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~1_combout ),
	.cout());
defparam \add_in_r_c~1 .lut_mask = 16'hAACC;
defparam \add_in_r_c~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~2 (
	.dataa(ram_in_reg_0_7),
	.datab(ram_in_reg_0_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~2_combout ),
	.cout());
defparam \add_in_r_d~2 .lut_mask = 16'hAACC;
defparam \add_in_r_d~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~2 (
	.dataa(ram_in_reg_0_5),
	.datab(ram_in_reg_0_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~2_combout ),
	.cout());
defparam \add_in_r_c~2 .lut_mask = 16'hAACC;
defparam \add_in_r_c~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~3 (
	.dataa(ram_in_reg_9_7),
	.datab(ram_in_reg_9_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~3_combout ),
	.cout());
defparam \add_in_r_d~3 .lut_mask = 16'hAACC;
defparam \add_in_r_d~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~3 (
	.dataa(ram_in_reg_9_5),
	.datab(ram_in_reg_9_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~3_combout ),
	.cout());
defparam \add_in_r_c~3 .lut_mask = 16'hAACC;
defparam \add_in_r_c~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~4 (
	.dataa(ram_in_reg_8_7),
	.datab(ram_in_reg_8_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~4_combout ),
	.cout());
defparam \add_in_r_d~4 .lut_mask = 16'hAACC;
defparam \add_in_r_d~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~4 (
	.dataa(ram_in_reg_8_5),
	.datab(ram_in_reg_8_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~4_combout ),
	.cout());
defparam \add_in_r_c~4 .lut_mask = 16'hAACC;
defparam \add_in_r_c~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~5 (
	.dataa(ram_in_reg_7_7),
	.datab(ram_in_reg_7_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~5_combout ),
	.cout());
defparam \add_in_r_d~5 .lut_mask = 16'hAACC;
defparam \add_in_r_d~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~5 (
	.dataa(ram_in_reg_7_5),
	.datab(ram_in_reg_7_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~5_combout ),
	.cout());
defparam \add_in_r_c~5 .lut_mask = 16'hAACC;
defparam \add_in_r_c~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~6 (
	.dataa(ram_in_reg_6_7),
	.datab(ram_in_reg_6_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~6_combout ),
	.cout());
defparam \add_in_r_d~6 .lut_mask = 16'hAACC;
defparam \add_in_r_d~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~6 (
	.dataa(ram_in_reg_6_5),
	.datab(ram_in_reg_6_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~6_combout ),
	.cout());
defparam \add_in_r_c~6 .lut_mask = 16'hAACC;
defparam \add_in_r_c~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~7 (
	.dataa(ram_in_reg_5_7),
	.datab(ram_in_reg_5_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~7_combout ),
	.cout());
defparam \add_in_r_d~7 .lut_mask = 16'hAACC;
defparam \add_in_r_d~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~7 (
	.dataa(ram_in_reg_5_5),
	.datab(ram_in_reg_5_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~7_combout ),
	.cout());
defparam \add_in_r_c~7 .lut_mask = 16'hAACC;
defparam \add_in_r_c~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~8 (
	.dataa(ram_in_reg_4_7),
	.datab(ram_in_reg_4_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~8_combout ),
	.cout());
defparam \add_in_r_d~8 .lut_mask = 16'hAACC;
defparam \add_in_r_d~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~8 (
	.dataa(ram_in_reg_4_5),
	.datab(ram_in_reg_4_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~8_combout ),
	.cout());
defparam \add_in_r_c~8 .lut_mask = 16'hAACC;
defparam \add_in_r_c~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_d~9 (
	.dataa(ram_in_reg_3_7),
	.datab(ram_in_reg_3_3),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_d~9_combout ),
	.cout());
defparam \add_in_r_d~9 .lut_mask = 16'hAACC;
defparam \add_in_r_d~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \add_in_r_c~9 (
	.dataa(ram_in_reg_3_5),
	.datab(ram_in_reg_3_1),
	.datac(gnd),
	.datad(\sign_sel[0]~q ),
	.cin(gnd),
	.combout(\add_in_r_c~9_combout ),
	.cout());
defparam \add_in_r_c~9 .lut_mask = 16'hAACC;
defparam \add_in_r_c~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \offset_counter[5]~28 (
	.dataa(tdl_arr_4),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\offset_counter[5]~28_combout ),
	.cout());
defparam \offset_counter[5]~28 .lut_mask = 16'hAAFF;
defparam \offset_counter[5]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\offset_counter[8]~q ),
	.datab(\offset_counter[9]~q ),
	.datac(\offset_counter[7]~q ),
	.datad(\offset_counter[0]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\offset_counter[4]~q ),
	.datab(\offset_counter[3]~q ),
	.datac(\offset_counter[2]~q ),
	.datad(\offset_counter[1]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFEFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\offset_counter[6]~q ),
	.datab(\offset_counter[5]~q ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFFFE;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_val_i~0 (
	.dataa(tdl_arr_4),
	.datab(\data_val_i~q ),
	.datac(gnd),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\data_val_i~0_combout ),
	.cout());
defparam \data_val_i~0 .lut_mask = 16'hEEFF;
defparam \data_val_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sign_vec[3]~1 (
	.dataa(\sign_sel[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sign_vec[3]~1_combout ),
	.cout());
defparam \sign_vec[3]~1 .lut_mask = 16'h5555;
defparam \sign_vec[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sign_vec[1]~2 (
	.dataa(\sign_sel[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sign_vec[1]~2_combout ),
	.cout());
defparam \sign_vec[1]~2 .lut_mask = 16'h5555;
defparam \sign_vec[1]~2 .sum_lutc_input = "datac";

dffeas \data_imag_o[0] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_0),
	.prn(vcc));
defparam \data_imag_o[0] .is_wysiwyg = "true";
defparam \data_imag_o[0] .power_up = "low";

dffeas \data_real_o[0] (
	.clk(clk),
	.d(\data_real_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_0),
	.prn(vcc));
defparam \data_real_o[0] .is_wysiwyg = "true";
defparam \data_real_o[0] .power_up = "low";

dffeas \data_imag_o[1] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_1),
	.prn(vcc));
defparam \data_imag_o[1] .is_wysiwyg = "true";
defparam \data_imag_o[1] .power_up = "low";

dffeas \data_real_o[1] (
	.clk(clk),
	.d(\data_real_o~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_1),
	.prn(vcc));
defparam \data_real_o[1] .is_wysiwyg = "true";
defparam \data_real_o[1] .power_up = "low";

dffeas \data_imag_o[2] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_2),
	.prn(vcc));
defparam \data_imag_o[2] .is_wysiwyg = "true";
defparam \data_imag_o[2] .power_up = "low";

dffeas \data_real_o[2] (
	.clk(clk),
	.d(\data_real_o~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_2),
	.prn(vcc));
defparam \data_real_o[2] .is_wysiwyg = "true";
defparam \data_real_o[2] .power_up = "low";

dffeas \data_imag_o[3] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_3),
	.prn(vcc));
defparam \data_imag_o[3] .is_wysiwyg = "true";
defparam \data_imag_o[3] .power_up = "low";

dffeas \data_real_o[3] (
	.clk(clk),
	.d(\data_real_o~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_3),
	.prn(vcc));
defparam \data_real_o[3] .is_wysiwyg = "true";
defparam \data_real_o[3] .power_up = "low";

dffeas \data_imag_o[4] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_4),
	.prn(vcc));
defparam \data_imag_o[4] .is_wysiwyg = "true";
defparam \data_imag_o[4] .power_up = "low";

dffeas \data_real_o[4] (
	.clk(clk),
	.d(\data_real_o~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_4),
	.prn(vcc));
defparam \data_real_o[4] .is_wysiwyg = "true";
defparam \data_real_o[4] .power_up = "low";

dffeas \data_imag_o[5] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_5),
	.prn(vcc));
defparam \data_imag_o[5] .is_wysiwyg = "true";
defparam \data_imag_o[5] .power_up = "low";

dffeas \data_real_o[5] (
	.clk(clk),
	.d(\data_real_o~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_5),
	.prn(vcc));
defparam \data_real_o[5] .is_wysiwyg = "true";
defparam \data_real_o[5] .power_up = "low";

dffeas \data_imag_o[6] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_6),
	.prn(vcc));
defparam \data_imag_o[6] .is_wysiwyg = "true";
defparam \data_imag_o[6] .power_up = "low";

dffeas \data_real_o[6] (
	.clk(clk),
	.d(\data_real_o~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_6),
	.prn(vcc));
defparam \data_real_o[6] .is_wysiwyg = "true";
defparam \data_real_o[6] .power_up = "low";

dffeas \data_imag_o[7] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_7),
	.prn(vcc));
defparam \data_imag_o[7] .is_wysiwyg = "true";
defparam \data_imag_o[7] .power_up = "low";

dffeas \data_real_o[7] (
	.clk(clk),
	.d(\data_real_o~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_7),
	.prn(vcc));
defparam \data_real_o[7] .is_wysiwyg = "true";
defparam \data_real_o[7] .power_up = "low";

dffeas \data_imag_o[8] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_8),
	.prn(vcc));
defparam \data_imag_o[8] .is_wysiwyg = "true";
defparam \data_imag_o[8] .power_up = "low";

dffeas \data_real_o[8] (
	.clk(clk),
	.d(\data_real_o~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_8),
	.prn(vcc));
defparam \data_real_o[8] .is_wysiwyg = "true";
defparam \data_real_o[8] .power_up = "low";

dffeas \data_imag_o[9] (
	.clk(clk),
	.d(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(data_imag_o_9),
	.prn(vcc));
defparam \data_imag_o[9] .is_wysiwyg = "true";
defparam \data_imag_o[9] .power_up = "low";

dffeas \data_real_o[9] (
	.clk(clk),
	.d(\data_real_o~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(data_real_o_9),
	.prn(vcc));
defparam \data_real_o[9] .is_wysiwyg = "true";
defparam \data_real_o[9] .power_up = "low";

cycloneive_lcell_comb \data_real_o~0 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~0_combout ),
	.cout());
defparam \data_real_o~0 .lut_mask = 16'hEEEE;
defparam \data_real_o~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~1 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~1_combout ),
	.cout());
defparam \data_real_o~1 .lut_mask = 16'hEEEE;
defparam \data_real_o~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~2 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~2_combout ),
	.cout());
defparam \data_real_o~2 .lut_mask = 16'hEEEE;
defparam \data_real_o~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~3 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~3_combout ),
	.cout());
defparam \data_real_o~3 .lut_mask = 16'hEEEE;
defparam \data_real_o~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~4 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~4_combout ),
	.cout());
defparam \data_real_o~4 .lut_mask = 16'hEEEE;
defparam \data_real_o~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~5 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~5_combout ),
	.cout());
defparam \data_real_o~5 .lut_mask = 16'hEEEE;
defparam \data_real_o~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~6 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~6_combout ),
	.cout());
defparam \data_real_o~6 .lut_mask = 16'hEEEE;
defparam \data_real_o~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~7 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~7_combout ),
	.cout());
defparam \data_real_o~7 .lut_mask = 16'hEEEE;
defparam \data_real_o~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~8 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~8_combout ),
	.cout());
defparam \data_real_o~8 .lut_mask = 16'hEEEE;
defparam \data_real_o~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_real_o~9 (
	.dataa(reset_n),
	.datab(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_real_o~9_combout ),
	.cout());
defparam \data_real_o~9 .lut_mask = 16'hEEEE;
defparam \data_real_o~9 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_pround_14 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_r_2,
	output_r_1,
	output_r_0,
	output_r_11,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_r_2;
input 	output_r_1;
input 	output_r_0;
input 	output_r_11;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_15 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.output_r_2(output_r_2),
	.output_r_1(output_r_1),
	.output_r_0(output_r_0),
	.output_r_11(output_r_11),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.output_r_8(output_r_8),
	.output_r_9(output_r_9),
	.output_r_10(output_r_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_15 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_r_2,
	output_r_1,
	output_r_0,
	output_r_11,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_r_2;
input 	output_r_1;
input 	output_r_0;
input 	output_r_11;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_8 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.output_r_2(output_r_2),
	.output_r_1(output_r_1),
	.output_r_0(output_r_0),
	.output_r_11(output_r_11),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.output_r_8(output_r_8),
	.output_r_9(output_r_9),
	.output_r_10(output_r_10),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_8 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_r_2,
	output_r_1,
	output_r_0,
	output_r_11,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_r_2;
input 	output_r_1;
input 	output_r_0;
input 	output_r_11;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(output_r_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(output_r_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(output_r_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(output_r_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(output_r_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(output_r_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(output_r_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(output_r_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(output_r_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(output_r_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(output_r_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(output_r_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(output_r_11),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_pround_15 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_i_2,
	output_i_1,
	output_i_0,
	output_i_11,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_10,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_i_2;
input 	output_i_1;
input 	output_i_0;
input 	output_i_11;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_10;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_LPM_ADD_SUB_16 \gbrnd:nev:gp:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.output_i_2(output_i_2),
	.output_i_1(output_i_1),
	.output_i_0(output_i_0),
	.output_i_11(output_i_11),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.output_i_8(output_i_8),
	.output_i_9(output_i_9),
	.output_i_10(output_i_10),
	.clken(global_clock_enable),
	.clock(clk));

endmodule

module fftsign_LPM_ADD_SUB_16 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_i_2,
	output_i_1,
	output_i_0,
	output_i_11,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_i_2;
input 	output_i_1;
input 	output_i_0;
input 	output_i_11;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_add_sub_inj_9 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.output_i_2(output_i_2),
	.output_i_1(output_i_1),
	.output_i_0(output_i_0),
	.output_i_11(output_i_11),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.output_i_8(output_i_8),
	.output_i_9(output_i_9),
	.output_i_10(output_i_10),
	.clken(clken),
	.clock(clock));

endmodule

module fftsign_add_sub_inj_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	output_i_2,
	output_i_1,
	output_i_0,
	output_i_11,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_10,
	clken,
	clock)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	output_i_2;
input 	output_i_1;
input 	output_i_0;
input 	output_i_11;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_10;
input 	clken;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ;
wire \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ;


dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(output_i_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h0055;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(output_i_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h005F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 (
	.dataa(output_i_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .lut_mask = 16'h00AF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 (
	.dataa(output_i_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15_cout ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 (
	.dataa(output_i_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~17 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 (
	.dataa(output_i_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~19 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 (
	.dataa(output_i_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~21 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 (
	.dataa(output_i_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~23 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 (
	.dataa(output_i_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~25 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 (
	.dataa(output_i_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~27 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 (
	.dataa(output_i_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~29 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .lut_mask = 16'h5AAF;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 (
	.dataa(output_i_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~31 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32_combout ),
	.cout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ));
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .lut_mask = 16'h5A5F;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 (
	.dataa(output_i_11),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~33 ),
	.combout(\fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34_combout ),
	.cout());
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .lut_mask = 16'h5A5A;
defparam \fft_ii_0|asj_fft_si_se_so_b_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~34 .sum_lutc_input = "cin";

endmodule

module fftsign_asj_fft_tdl_bit_1 (
	data_in,
	global_clock_enable,
	tdl_arr_4,
	clk)/* synthesis synthesis_greybox=1 */;
input 	data_in;
input 	global_clock_enable;
output 	tdl_arr_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

endmodule

module fftsign_asj_fft_lpprdadgen (
	lpp_c_i,
	global_clock_enable,
	tdl_arr_4,
	tdl_arr_0_4,
	tdl_arr_1_4,
	en_d1,
	rd_addr_d_0,
	rd_addr_d_1,
	rd_addr_d_2,
	rd_addr_d_3,
	rd_addr_d_4,
	rd_addr_d_5,
	sw_0,
	sw_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	lpp_c_i;
input 	global_clock_enable;
output 	tdl_arr_4;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
output 	en_d1;
output 	rd_addr_d_0;
output 	rd_addr_d_1;
output 	rd_addr_d_2;
output 	rd_addr_d_3;
output 	rd_addr_d_4;
output 	rd_addr_d_5;
output 	sw_0;
output 	sw_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \en_d~0_combout ;
wire \count[0]~8_combout ;
wire \en_i~0_combout ;
wire \en_i~q ;
wire \counter~0_combout ;
wire \count[0]~q ;
wire \count[0]~9 ;
wire \count[1]~10_combout ;
wire \count[1]~q ;
wire \count[1]~11 ;
wire \count[2]~12_combout ;
wire \count[2]~q ;
wire \count[2]~13 ;
wire \count[3]~14_combout ;
wire \count[3]~q ;
wire \count[3]~15 ;
wire \count[4]~16_combout ;
wire \count[4]~q ;
wire \count[4]~17 ;
wire \count[5]~18_combout ;
wire \count[5]~q ;
wire \count[5]~19 ;
wire \count[6]~20_combout ;
wire \count[6]~q ;
wire \count[6]~21 ;
wire \count[7]~22_combout ;
wire \count[7]~q ;
wire \Add3~0_combout ;
wire \Add3~1_combout ;
wire \Add3~2_combout ;
wire \Add3~3_combout ;


fftsign_asj_fft_tdl_rst \gen_M4K:delay_swd (
	.global_clock_enable(global_clock_enable),
	.tdl_arr_0_4(tdl_arr_0_4),
	.tdl_arr_1_4(tdl_arr_1_4),
	.sw_0(sw_0),
	.sw_1(sw_1),
	.clk(clk),
	.reset_n(reset_n));

fftsign_asj_fft_tdl_bit_rst_4 delay_en(
	.en_i(\en_i~q ),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_4(tdl_arr_4),
	.clk(clk),
	.reset_n(reset_n));

dffeas en_d(
	.clk(clk),
	.d(\en_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(en_d1),
	.prn(vcc));
defparam en_d.is_wysiwyg = "true";
defparam en_d.power_up = "low";

dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

dffeas \rd_addr_d[2] (
	.clk(clk),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_2),
	.prn(vcc));
defparam \rd_addr_d[2] .is_wysiwyg = "true";
defparam \rd_addr_d[2] .power_up = "low";

dffeas \rd_addr_d[3] (
	.clk(clk),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_3),
	.prn(vcc));
defparam \rd_addr_d[3] .is_wysiwyg = "true";
defparam \rd_addr_d[3] .power_up = "low";

dffeas \rd_addr_d[4] (
	.clk(clk),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_4),
	.prn(vcc));
defparam \rd_addr_d[4] .is_wysiwyg = "true";
defparam \rd_addr_d[4] .power_up = "low";

dffeas \rd_addr_d[5] (
	.clk(clk),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rd_addr_d_5),
	.prn(vcc));
defparam \rd_addr_d[5] .is_wysiwyg = "true";
defparam \rd_addr_d[5] .power_up = "low";

dffeas \sw[0] (
	.clk(clk),
	.d(\Add3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \sw[1] (
	.clk(clk),
	.d(\Add3~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(sw_1),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

cycloneive_lcell_comb \en_d~0 (
	.dataa(reset_n),
	.datab(lpp_c_i),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\en_d~0_combout ),
	.cout());
defparam \en_d~0 .lut_mask = 16'hEEEE;
defparam \en_d~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~8 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~8_combout ),
	.cout(\count[0]~9 ));
defparam \count[0]~8 .lut_mask = 16'h55AA;
defparam \count[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \en_i~0 (
	.dataa(lpp_c_i),
	.datab(gnd),
	.datac(gnd),
	.datad(en_d1),
	.cin(gnd),
	.combout(\en_i~0_combout ),
	.cout());
defparam \en_i~0 .lut_mask = 16'hAAFF;
defparam \en_i~0 .sum_lutc_input = "datac";

dffeas en_i(
	.clk(clk),
	.d(\en_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\en_i~q ),
	.prn(vcc));
defparam en_i.is_wysiwyg = "true";
defparam en_i.power_up = "low";

cycloneive_lcell_comb \counter~0 (
	.dataa(\en_i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\counter~0_combout ),
	.cout());
defparam \counter~0 .lut_mask = 16'hAAFF;
defparam \counter~0 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \count[1]~10 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~9 ),
	.combout(\count[1]~10_combout ),
	.cout(\count[1]~11 ));
defparam \count[1]~10 .lut_mask = 16'h5A5F;
defparam \count[1]~10 .sum_lutc_input = "cin";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \count[2]~12 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~11 ),
	.combout(\count[2]~12_combout ),
	.cout(\count[2]~13 ));
defparam \count[2]~12 .lut_mask = 16'h5AAF;
defparam \count[2]~12 .sum_lutc_input = "cin";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count[3]~14 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~13 ),
	.combout(\count[3]~14_combout ),
	.cout(\count[3]~15 ));
defparam \count[3]~14 .lut_mask = 16'h5A5F;
defparam \count[3]~14 .sum_lutc_input = "cin";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count[4]~16 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~15 ),
	.combout(\count[4]~16_combout ),
	.cout(\count[4]~17 ));
defparam \count[4]~16 .lut_mask = 16'h5AAF;
defparam \count[4]~16 .sum_lutc_input = "cin";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count[5]~18 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~17 ),
	.combout(\count[5]~18_combout ),
	.cout(\count[5]~19 ));
defparam \count[5]~18 .lut_mask = 16'h5A5F;
defparam \count[5]~18 .sum_lutc_input = "cin";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count[6]~20 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~19 ),
	.combout(\count[6]~20_combout ),
	.cout(\count[6]~21 ));
defparam \count[6]~20 .lut_mask = 16'h5AAF;
defparam \count[6]~20 .sum_lutc_input = "cin";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count[7]~22 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[6]~21 ),
	.combout(\count[7]~22_combout ),
	.cout());
defparam \count[7]~22 .lut_mask = 16'h5A5A;
defparam \count[7]~22 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter~0_combout ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \Add3~0 (
	.dataa(\count[2]~q ),
	.datab(\count[4]~q ),
	.datac(\count[6]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h6996;
defparam \Add3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~1 (
	.dataa(\count[2]~q ),
	.datab(\count[4]~q ),
	.datac(\count[6]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'h6996;
defparam \Add3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~2 (
	.dataa(\count[3]~q ),
	.datab(\count[5]~q ),
	.datac(\count[7]~q ),
	.datad(\count[1]~q ),
	.cin(gnd),
	.combout(\Add3~2_combout ),
	.cout());
defparam \Add3~2 .lut_mask = 16'h6996;
defparam \Add3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add3~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Add3~1_combout ),
	.datad(\Add3~2_combout ),
	.cin(gnd),
	.combout(\Add3~3_combout ),
	.cout());
defparam \Add3~3 .lut_mask = 16'h0FF0;
defparam \Add3~3 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_rst_4 (
	en_i,
	global_clock_enable,
	tdl_arr_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	en_i;
input 	global_clock_enable;
output 	tdl_arr_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~4_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(en_i),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_rst (
	global_clock_enable,
	tdl_arr_0_4,
	tdl_arr_1_4,
	sw_0,
	sw_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
input 	sw_0;
input 	sw_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~8_combout ;
wire \tdl_arr[0][0]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[1][0]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[2][0]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[3][0]~q ;
wire \tdl_arr~0_combout ;
wire \tdl_arr~9_combout ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[1][1]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[2][1]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[3][1]~q ;
wire \tdl_arr~1_combout ;


dffeas \tdl_arr[4][0] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0_4),
	.prn(vcc));
defparam \tdl_arr[4][0] .is_wysiwyg = "true";
defparam \tdl_arr[4][0] .power_up = "low";

dffeas \tdl_arr[4][1] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_1_4),
	.prn(vcc));
defparam \tdl_arr[4][1] .is_wysiwyg = "true";
defparam \tdl_arr[4][1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(sw_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][0]~q ),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[2][0] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][0]~q ),
	.prn(vcc));
defparam \tdl_arr[2][0] .is_wysiwyg = "true";
defparam \tdl_arr[2][0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[3][0] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][0]~q ),
	.prn(vcc));
defparam \tdl_arr[3][0] .is_wysiwyg = "true";
defparam \tdl_arr[3][0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(sw_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1][1]~q ),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[2][1] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2][1]~q ),
	.prn(vcc));
defparam \tdl_arr[2][1] .is_wysiwyg = "true";
defparam \tdl_arr[2][1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[3][1] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3][1]~q ),
	.prn(vcc));
defparam \tdl_arr[3][1] .is_wysiwyg = "true";
defparam \tdl_arr[3][1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_m_k_counter (
	rdy_for_next_block,
	blk_done_int1,
	global_clock_enable,
	tdl_arr_0,
	p_2,
	p_0,
	p_1,
	k_count_4,
	k_count_0,
	k_count_2,
	k_count_6,
	k_count_1,
	k_count_3,
	k_count_5,
	k_count_7,
	data_rdy_vec_4,
	next_pass_i1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	rdy_for_next_block;
output 	blk_done_int1;
input 	global_clock_enable;
input 	tdl_arr_0;
output 	p_2;
output 	p_0;
output 	p_1;
output 	k_count_4;
output 	k_count_0;
output 	k_count_2;
output 	k_count_6;
output 	k_count_1;
output 	k_count_3;
output 	k_count_5;
output 	k_count_7;
input 	data_rdy_vec_4;
output 	next_pass_i1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \k[0]~8_combout ;
wire \next_block_d2~q ;
wire \next_block_d3~q ;
wire \next_block_d4~q ;
wire \cnt_k~0_combout ;
wire \cnt_k~1_combout ;
wire \next_pass_id~0_combout ;
wire \del_npi_cnt[0]~6_combout ;
wire \del_npi_cnt[0]~q ;
wire \del_npi_cnt[0]~7 ;
wire \del_npi_cnt[1]~8_combout ;
wire \del_npi_cnt[1]~q ;
wire \del_npi_cnt[1]~9 ;
wire \del_npi_cnt[2]~10_combout ;
wire \del_npi_cnt[2]~q ;
wire \del_npi_cnt[2]~11 ;
wire \del_npi_cnt[3]~12_combout ;
wire \del_npi_cnt[3]~q ;
wire \next_pass_id~1_combout ;
wire \del_npi_cnt[3]~13 ;
wire \del_npi_cnt[4]~14_combout ;
wire \del_npi_cnt[4]~q ;
wire \next_pass_id~2_combout ;
wire \next_pass_id~q ;
wire \Selector2~0_combout ;
wire \k_state.HOLD~q ;
wire \k_state.IDLE~0_combout ;
wire \k_state.IDLE~1_combout ;
wire \k_state.IDLE~q ;
wire \k[0]~20_combout ;
wire \k[0]~q ;
wire \k[0]~9 ;
wire \k[1]~10_combout ;
wire \k[1]~q ;
wire \k[1]~11 ;
wire \k[2]~12_combout ;
wire \k[2]~q ;
wire \k[2]~13 ;
wire \k[3]~14_combout ;
wire \k[3]~q ;
wire \k[3]~15 ;
wire \k[4]~16_combout ;
wire \k[4]~q ;
wire \k[4]~17 ;
wire \k[5]~18_combout ;
wire \k[5]~q ;
wire \Equal3~0_combout ;
wire \k[5]~19 ;
wire \k[6]~21_combout ;
wire \k[6]~q ;
wire \k[6]~22 ;
wire \k[7]~23_combout ;
wire \k[7]~q ;
wire \Equal3~1_combout ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \k_state.RUN_CNT~q ;
wire \k_state~8_combout ;
wire \k_state.NEXT_PASS_UPD~q ;
wire \blk_done_int~0_combout ;
wire \p~2_combout ;
wire \p~3_combout ;
wire \p[2]~4_combout ;
wire \p~5_combout ;
wire \p~6_combout ;
wire \p~7_combout ;
wire \next_pass_i~0_combout ;


dffeas blk_done_int(
	.clk(clk),
	.d(\blk_done_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(blk_done_int1),
	.prn(vcc));
defparam blk_done_int.is_wysiwyg = "true";
defparam blk_done_int.power_up = "low";

dffeas \p[2] (
	.clk(clk),
	.d(\p~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[2]~4_combout ),
	.q(p_2),
	.prn(vcc));
defparam \p[2] .is_wysiwyg = "true";
defparam \p[2] .power_up = "low";

dffeas \p[0] (
	.clk(clk),
	.d(\p~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[2]~4_combout ),
	.q(p_0),
	.prn(vcc));
defparam \p[0] .is_wysiwyg = "true";
defparam \p[0] .power_up = "low";

dffeas \p[1] (
	.clk(clk),
	.d(\p~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[2]~4_combout ),
	.q(p_1),
	.prn(vcc));
defparam \p[1] .is_wysiwyg = "true";
defparam \p[1] .power_up = "low";

dffeas \k_count[4] (
	.clk(clk),
	.d(\k[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_4),
	.prn(vcc));
defparam \k_count[4] .is_wysiwyg = "true";
defparam \k_count[4] .power_up = "low";

dffeas \k_count[0] (
	.clk(clk),
	.d(\k[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_0),
	.prn(vcc));
defparam \k_count[0] .is_wysiwyg = "true";
defparam \k_count[0] .power_up = "low";

dffeas \k_count[2] (
	.clk(clk),
	.d(\k[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_2),
	.prn(vcc));
defparam \k_count[2] .is_wysiwyg = "true";
defparam \k_count[2] .power_up = "low";

dffeas \k_count[6] (
	.clk(clk),
	.d(\k[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_6),
	.prn(vcc));
defparam \k_count[6] .is_wysiwyg = "true";
defparam \k_count[6] .power_up = "low";

dffeas \k_count[1] (
	.clk(clk),
	.d(\k[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_1),
	.prn(vcc));
defparam \k_count[1] .is_wysiwyg = "true";
defparam \k_count[1] .power_up = "low";

dffeas \k_count[3] (
	.clk(clk),
	.d(\k[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_3),
	.prn(vcc));
defparam \k_count[3] .is_wysiwyg = "true";
defparam \k_count[3] .power_up = "low";

dffeas \k_count[5] (
	.clk(clk),
	.d(\k[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_5),
	.prn(vcc));
defparam \k_count[5] .is_wysiwyg = "true";
defparam \k_count[5] .power_up = "low";

dffeas \k_count[7] (
	.clk(clk),
	.d(\k[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(k_count_7),
	.prn(vcc));
defparam \k_count[7] .is_wysiwyg = "true";
defparam \k_count[7] .power_up = "low";

dffeas next_pass_i(
	.clk(clk),
	.d(\next_pass_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(next_pass_i1),
	.prn(vcc));
defparam next_pass_i.is_wysiwyg = "true";
defparam next_pass_i.power_up = "low";

cycloneive_lcell_comb \k[0]~8 (
	.dataa(\k[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\k[0]~8_combout ),
	.cout(\k[0]~9 ));
defparam \k[0]~8 .lut_mask = 16'h55AA;
defparam \k[0]~8 .sum_lutc_input = "datac";

dffeas next_block_d2(
	.clk(clk),
	.d(tdl_arr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_block_d2~q ),
	.prn(vcc));
defparam next_block_d2.is_wysiwyg = "true";
defparam next_block_d2.power_up = "low";

dffeas next_block_d3(
	.clk(clk),
	.d(\next_block_d2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_block_d3~q ),
	.prn(vcc));
defparam next_block_d3.is_wysiwyg = "true";
defparam next_block_d3.power_up = "low";

dffeas next_block_d4(
	.clk(clk),
	.d(\next_block_d3~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_block_d4~q ),
	.prn(vcc));
defparam next_block_d4.is_wysiwyg = "true";
defparam next_block_d4.power_up = "low";

cycloneive_lcell_comb \cnt_k~0 (
	.dataa(rdy_for_next_block),
	.datab(\next_block_d4~q ),
	.datac(\next_block_d3~q ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\cnt_k~0_combout ),
	.cout());
defparam \cnt_k~0 .lut_mask = 16'hFEFF;
defparam \cnt_k~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cnt_k~1 (
	.dataa(tdl_arr_0),
	.datab(\cnt_k~0_combout ),
	.datac(\next_block_d2~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\cnt_k~1_combout ),
	.cout());
defparam \cnt_k~1 .lut_mask = 16'hFEFE;
defparam \cnt_k~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_pass_id~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\next_pass_id~0_combout ),
	.cout());
defparam \next_pass_id~0 .lut_mask = 16'hFFFE;
defparam \next_pass_id~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_npi_cnt[0]~6 (
	.dataa(\del_npi_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\del_npi_cnt[0]~6_combout ),
	.cout(\del_npi_cnt[0]~7 ));
defparam \del_npi_cnt[0]~6 .lut_mask = 16'h55AA;
defparam \del_npi_cnt[0]~6 .sum_lutc_input = "datac";

dffeas \del_npi_cnt[0] (
	.clk(clk),
	.d(\del_npi_cnt[0]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[0]~q ),
	.prn(vcc));
defparam \del_npi_cnt[0] .is_wysiwyg = "true";
defparam \del_npi_cnt[0] .power_up = "low";

cycloneive_lcell_comb \del_npi_cnt[1]~8 (
	.dataa(\del_npi_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[0]~7 ),
	.combout(\del_npi_cnt[1]~8_combout ),
	.cout(\del_npi_cnt[1]~9 ));
defparam \del_npi_cnt[1]~8 .lut_mask = 16'h5A5F;
defparam \del_npi_cnt[1]~8 .sum_lutc_input = "cin";

dffeas \del_npi_cnt[1] (
	.clk(clk),
	.d(\del_npi_cnt[1]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[1]~q ),
	.prn(vcc));
defparam \del_npi_cnt[1] .is_wysiwyg = "true";
defparam \del_npi_cnt[1] .power_up = "low";

cycloneive_lcell_comb \del_npi_cnt[2]~10 (
	.dataa(\del_npi_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[1]~9 ),
	.combout(\del_npi_cnt[2]~10_combout ),
	.cout(\del_npi_cnt[2]~11 ));
defparam \del_npi_cnt[2]~10 .lut_mask = 16'h5AAF;
defparam \del_npi_cnt[2]~10 .sum_lutc_input = "cin";

dffeas \del_npi_cnt[2] (
	.clk(clk),
	.d(\del_npi_cnt[2]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[2]~q ),
	.prn(vcc));
defparam \del_npi_cnt[2] .is_wysiwyg = "true";
defparam \del_npi_cnt[2] .power_up = "low";

cycloneive_lcell_comb \del_npi_cnt[3]~12 (
	.dataa(\del_npi_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\del_npi_cnt[2]~11 ),
	.combout(\del_npi_cnt[3]~12_combout ),
	.cout(\del_npi_cnt[3]~13 ));
defparam \del_npi_cnt[3]~12 .lut_mask = 16'h5A5F;
defparam \del_npi_cnt[3]~12 .sum_lutc_input = "cin";

dffeas \del_npi_cnt[3] (
	.clk(clk),
	.d(\del_npi_cnt[3]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[3]~q ),
	.prn(vcc));
defparam \del_npi_cnt[3] .is_wysiwyg = "true";
defparam \del_npi_cnt[3] .power_up = "low";

cycloneive_lcell_comb \next_pass_id~1 (
	.dataa(\del_npi_cnt[0]~q ),
	.datab(\del_npi_cnt[1]~q ),
	.datac(\del_npi_cnt[3]~q ),
	.datad(\del_npi_cnt[2]~q ),
	.cin(gnd),
	.combout(\next_pass_id~1_combout ),
	.cout());
defparam \next_pass_id~1 .lut_mask = 16'hFEFF;
defparam \next_pass_id~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \del_npi_cnt[4]~14 (
	.dataa(\del_npi_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\del_npi_cnt[3]~13 ),
	.combout(\del_npi_cnt[4]~14_combout ),
	.cout());
defparam \del_npi_cnt[4]~14 .lut_mask = 16'h5A5A;
defparam \del_npi_cnt[4]~14 .sum_lutc_input = "cin";

dffeas \del_npi_cnt[4] (
	.clk(clk),
	.d(\del_npi_cnt[4]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\k_state.HOLD~q ),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\del_npi_cnt[4]~q ),
	.prn(vcc));
defparam \del_npi_cnt[4] .is_wysiwyg = "true";
defparam \del_npi_cnt[4] .power_up = "low";

cycloneive_lcell_comb \next_pass_id~2 (
	.dataa(\next_pass_id~0_combout ),
	.datab(\next_pass_id~1_combout ),
	.datac(gnd),
	.datad(\del_npi_cnt[4]~q ),
	.cin(gnd),
	.combout(\next_pass_id~2_combout ),
	.cout());
defparam \next_pass_id~2 .lut_mask = 16'hEEFF;
defparam \next_pass_id~2 .sum_lutc_input = "datac";

dffeas next_pass_id(
	.clk(clk),
	.d(\next_pass_id~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\next_pass_id~q ),
	.prn(vcc));
defparam next_pass_id.is_wysiwyg = "true";
defparam next_pass_id.power_up = "low";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\k_state.NEXT_PASS_UPD~q ),
	.datab(data_rdy_vec_4),
	.datac(\k_state.HOLD~q ),
	.datad(\next_pass_id~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \k_state.HOLD (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.HOLD~q ),
	.prn(vcc));
defparam \k_state.HOLD .is_wysiwyg = "true";
defparam \k_state.HOLD .power_up = "low";

cycloneive_lcell_comb \k_state.IDLE~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(\next_pass_id~q ),
	.datac(\k_state.IDLE~q ),
	.datad(data_rdy_vec_4),
	.cin(gnd),
	.combout(\k_state.IDLE~0_combout ),
	.cout());
defparam \k_state.IDLE~0 .lut_mask = 16'hBFFF;
defparam \k_state.IDLE~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k_state.IDLE~1 (
	.dataa(\k_state.IDLE~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\k_state.IDLE~1_combout ),
	.cout());
defparam \k_state.IDLE~1 .lut_mask = 16'hFF55;
defparam \k_state.IDLE~1 .sum_lutc_input = "datac";

dffeas \k_state.IDLE (
	.clk(clk),
	.d(\k_state.IDLE~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.IDLE~q ),
	.prn(vcc));
defparam \k_state.IDLE .is_wysiwyg = "true";
defparam \k_state.IDLE .power_up = "low";

cycloneive_lcell_comb \k[0]~20 (
	.dataa(global_clock_enable),
	.datab(\k_state.HOLD~q ),
	.datac(\k_state.IDLE~q ),
	.datad(\cnt_k~1_combout ),
	.cin(gnd),
	.combout(\k[0]~20_combout ),
	.cout());
defparam \k[0]~20 .lut_mask = 16'hFFFB;
defparam \k[0]~20 .sum_lutc_input = "datac";

dffeas \k[0] (
	.clk(clk),
	.d(\k[0]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[0]~q ),
	.prn(vcc));
defparam \k[0] .is_wysiwyg = "true";
defparam \k[0] .power_up = "low";

cycloneive_lcell_comb \k[1]~10 (
	.dataa(\k[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[0]~9 ),
	.combout(\k[1]~10_combout ),
	.cout(\k[1]~11 ));
defparam \k[1]~10 .lut_mask = 16'h5A5F;
defparam \k[1]~10 .sum_lutc_input = "cin";

dffeas \k[1] (
	.clk(clk),
	.d(\k[1]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[1]~q ),
	.prn(vcc));
defparam \k[1] .is_wysiwyg = "true";
defparam \k[1] .power_up = "low";

cycloneive_lcell_comb \k[2]~12 (
	.dataa(\k[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[1]~11 ),
	.combout(\k[2]~12_combout ),
	.cout(\k[2]~13 ));
defparam \k[2]~12 .lut_mask = 16'h5AAF;
defparam \k[2]~12 .sum_lutc_input = "cin";

dffeas \k[2] (
	.clk(clk),
	.d(\k[2]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[2]~q ),
	.prn(vcc));
defparam \k[2] .is_wysiwyg = "true";
defparam \k[2] .power_up = "low";

cycloneive_lcell_comb \k[3]~14 (
	.dataa(\k[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[2]~13 ),
	.combout(\k[3]~14_combout ),
	.cout(\k[3]~15 ));
defparam \k[3]~14 .lut_mask = 16'h5A5F;
defparam \k[3]~14 .sum_lutc_input = "cin";

dffeas \k[3] (
	.clk(clk),
	.d(\k[3]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[3]~q ),
	.prn(vcc));
defparam \k[3] .is_wysiwyg = "true";
defparam \k[3] .power_up = "low";

cycloneive_lcell_comb \k[4]~16 (
	.dataa(\k[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[3]~15 ),
	.combout(\k[4]~16_combout ),
	.cout(\k[4]~17 ));
defparam \k[4]~16 .lut_mask = 16'h5AAF;
defparam \k[4]~16 .sum_lutc_input = "cin";

dffeas \k[4] (
	.clk(clk),
	.d(\k[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[4]~q ),
	.prn(vcc));
defparam \k[4] .is_wysiwyg = "true";
defparam \k[4] .power_up = "low";

cycloneive_lcell_comb \k[5]~18 (
	.dataa(\k[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[4]~17 ),
	.combout(\k[5]~18_combout ),
	.cout(\k[5]~19 ));
defparam \k[5]~18 .lut_mask = 16'h5A5F;
defparam \k[5]~18 .sum_lutc_input = "cin";

dffeas \k[5] (
	.clk(clk),
	.d(\k[5]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[5]~q ),
	.prn(vcc));
defparam \k[5] .is_wysiwyg = "true";
defparam \k[5] .power_up = "low";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(\k[5]~q ),
	.datab(\k[1]~q ),
	.datac(\k[3]~q ),
	.datad(\k[0]~q ),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hFEFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \k[6]~21 (
	.dataa(\k[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\k[5]~19 ),
	.combout(\k[6]~21_combout ),
	.cout(\k[6]~22 ));
defparam \k[6]~21 .lut_mask = 16'h5AAF;
defparam \k[6]~21 .sum_lutc_input = "cin";

dffeas \k[6] (
	.clk(clk),
	.d(\k[6]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[6]~q ),
	.prn(vcc));
defparam \k[6] .is_wysiwyg = "true";
defparam \k[6] .power_up = "low";

cycloneive_lcell_comb \k[7]~23 (
	.dataa(\k[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\k[6]~22 ),
	.combout(\k[7]~23_combout ),
	.cout());
defparam \k[7]~23 .lut_mask = 16'h5A5A;
defparam \k[7]~23 .sum_lutc_input = "cin";

dffeas \k[7] (
	.clk(clk),
	.d(\k[7]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\cnt_k~1_combout ),
	.sload(gnd),
	.ena(\k[0]~20_combout ),
	.q(\k[7]~q ),
	.prn(vcc));
defparam \k[7] .is_wysiwyg = "true";
defparam \k[7] .power_up = "low";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(\k[2]~q ),
	.datab(\k[4]~q ),
	.datac(\k[7]~q ),
	.datad(\k[6]~q ),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
defparam \Equal3~1 .lut_mask = 16'hFFFE;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\k_state.HOLD~q ),
	.datab(\next_pass_id~q ),
	.datac(data_rdy_vec_4),
	.datad(\k_state.IDLE~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\Selector1~0_combout ),
	.datab(\k_state.RUN_CNT~q ),
	.datac(\Equal3~0_combout ),
	.datad(\Equal3~1_combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

dffeas \k_state.RUN_CNT (
	.clk(clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.RUN_CNT~q ),
	.prn(vcc));
defparam \k_state.RUN_CNT .is_wysiwyg = "true";
defparam \k_state.RUN_CNT .power_up = "low";

cycloneive_lcell_comb \k_state~8 (
	.dataa(reset_n),
	.datab(\Equal3~0_combout ),
	.datac(\Equal3~1_combout ),
	.datad(\k_state.RUN_CNT~q ),
	.cin(gnd),
	.combout(\k_state~8_combout ),
	.cout());
defparam \k_state~8 .lut_mask = 16'hFFFE;
defparam \k_state~8 .sum_lutc_input = "datac";

dffeas \k_state.NEXT_PASS_UPD (
	.clk(clk),
	.d(\k_state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\k_state.NEXT_PASS_UPD~q ),
	.prn(vcc));
defparam \k_state.NEXT_PASS_UPD .is_wysiwyg = "true";
defparam \k_state.NEXT_PASS_UPD .power_up = "low";

cycloneive_lcell_comb \blk_done_int~0 (
	.dataa(p_2),
	.datab(\k_state.NEXT_PASS_UPD~q ),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\blk_done_int~0_combout ),
	.cout());
defparam \blk_done_int~0 .lut_mask = 16'hEFFF;
defparam \blk_done_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~2 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(rdy_for_next_block),
	.cin(gnd),
	.combout(\p~2_combout ),
	.cout());
defparam \p~2 .lut_mask = 16'hAAFF;
defparam \p~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~3 (
	.dataa(\p~2_combout ),
	.datab(p_2),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\p~3_combout ),
	.cout());
defparam \p~3 .lut_mask = 16'hEBBE;
defparam \p~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p[2]~4 (
	.dataa(global_clock_enable),
	.datab(\p~2_combout ),
	.datac(data_rdy_vec_4),
	.datad(next_pass_i1),
	.cin(gnd),
	.combout(\p[2]~4_combout ),
	.cout());
defparam \p[2]~4 .lut_mask = 16'hFFFB;
defparam \p[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~5 (
	.dataa(rdy_for_next_block),
	.datab(p_1),
	.datac(p_2),
	.datad(p_0),
	.cin(gnd),
	.combout(\p~5_combout ),
	.cout());
defparam \p~5 .lut_mask = 16'hEFFF;
defparam \p~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~6 (
	.dataa(reset_n),
	.datab(\p~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p~6_combout ),
	.cout());
defparam \p~6 .lut_mask = 16'hEEEE;
defparam \p~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \p~7 (
	.dataa(reset_n),
	.datab(rdy_for_next_block),
	.datac(p_0),
	.datad(p_1),
	.cin(gnd),
	.combout(\p~7_combout ),
	.cout());
defparam \p~7 .lut_mask = 16'hBFFB;
defparam \p~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_pass_i~0 (
	.dataa(reset_n),
	.datab(\k_state.NEXT_PASS_UPD~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pass_i~0_combout ),
	.cout());
defparam \next_pass_i~0 .lut_mask = 16'hEEEE;
defparam \next_pass_i~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_2 (
	data_in,
	global_clock_enable,
	tdl_arr_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	data_in;
input 	global_clock_enable;
output 	tdl_arr_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module fftsign_asj_fft_tdl_bit_3 (
	data_in,
	global_clock_enable,
	tdl_arr_23,
	clk)/* synthesis synthesis_greybox=1 */;
input 	data_in;
input 	global_clock_enable;
output 	tdl_arr_23;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;
wire \tdl_arr[8]~q ;
wire \tdl_arr[9]~q ;
wire \tdl_arr[10]~q ;
wire \tdl_arr[11]~q ;
wire \tdl_arr[12]~q ;
wire \tdl_arr[13]~q ;
wire \tdl_arr[14]~q ;
wire \tdl_arr[15]~q ;
wire \tdl_arr[16]~q ;
wire \tdl_arr[17]~q ;
wire \tdl_arr[18]~q ;
wire \tdl_arr[19]~q ;
wire \tdl_arr[20]~q ;
wire \tdl_arr[21]~q ;
wire \tdl_arr[22]~q ;


dffeas \tdl_arr[23] (
	.clk(clk),
	.d(\tdl_arr[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_23),
	.prn(vcc));
defparam \tdl_arr[23] .is_wysiwyg = "true";
defparam \tdl_arr[23] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(data_in),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[11]~q ),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

dffeas \tdl_arr[12] (
	.clk(clk),
	.d(\tdl_arr[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[12]~q ),
	.prn(vcc));
defparam \tdl_arr[12] .is_wysiwyg = "true";
defparam \tdl_arr[12] .power_up = "low";

dffeas \tdl_arr[13] (
	.clk(clk),
	.d(\tdl_arr[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[13]~q ),
	.prn(vcc));
defparam \tdl_arr[13] .is_wysiwyg = "true";
defparam \tdl_arr[13] .power_up = "low";

dffeas \tdl_arr[14] (
	.clk(clk),
	.d(\tdl_arr[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[14]~q ),
	.prn(vcc));
defparam \tdl_arr[14] .is_wysiwyg = "true";
defparam \tdl_arr[14] .power_up = "low";

dffeas \tdl_arr[15] (
	.clk(clk),
	.d(\tdl_arr[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[15]~q ),
	.prn(vcc));
defparam \tdl_arr[15] .is_wysiwyg = "true";
defparam \tdl_arr[15] .power_up = "low";

dffeas \tdl_arr[16] (
	.clk(clk),
	.d(\tdl_arr[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[16]~q ),
	.prn(vcc));
defparam \tdl_arr[16] .is_wysiwyg = "true";
defparam \tdl_arr[16] .power_up = "low";

dffeas \tdl_arr[17] (
	.clk(clk),
	.d(\tdl_arr[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[17]~q ),
	.prn(vcc));
defparam \tdl_arr[17] .is_wysiwyg = "true";
defparam \tdl_arr[17] .power_up = "low";

dffeas \tdl_arr[18] (
	.clk(clk),
	.d(\tdl_arr[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[18]~q ),
	.prn(vcc));
defparam \tdl_arr[18] .is_wysiwyg = "true";
defparam \tdl_arr[18] .power_up = "low";

dffeas \tdl_arr[19] (
	.clk(clk),
	.d(\tdl_arr[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[19]~q ),
	.prn(vcc));
defparam \tdl_arr[19] .is_wysiwyg = "true";
defparam \tdl_arr[19] .power_up = "low";

dffeas \tdl_arr[20] (
	.clk(clk),
	.d(\tdl_arr[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[20]~q ),
	.prn(vcc));
defparam \tdl_arr[20] .is_wysiwyg = "true";
defparam \tdl_arr[20] .power_up = "low";

dffeas \tdl_arr[21] (
	.clk(clk),
	.d(\tdl_arr[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[21]~q ),
	.prn(vcc));
defparam \tdl_arr[21] .is_wysiwyg = "true";
defparam \tdl_arr[21] .power_up = "low";

dffeas \tdl_arr[22] (
	.clk(clk),
	.d(\tdl_arr[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[22]~q ),
	.prn(vcc));
defparam \tdl_arr[22] .is_wysiwyg = "true";
defparam \tdl_arr[22] .power_up = "low";

endmodule

module fftsign_asj_fft_tdl_bit_rst_5 (
	global_clock_enable,
	tdl_arr_9,
	next_pass_i,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_9;
input 	next_pass_i;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~9_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~8_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~7_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~6_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[6]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[7]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[8]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_9),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~9 (
	.dataa(reset_n),
	.datab(next_pass_i),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~9_combout ),
	.cout());
defparam \tdl_arr~9 .lut_mask = 16'hEEEE;
defparam \tdl_arr~9 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~8 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~8_combout ),
	.cout());
defparam \tdl_arr~8 .lut_mask = 16'hEEEE;
defparam \tdl_arr~8 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~7 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~7_combout ),
	.cout());
defparam \tdl_arr~7 .lut_mask = 16'hEEEE;
defparam \tdl_arr~7 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_tdl_bit_rst_6 (
	global_clock_enable,
	tdl_arr_4,
	tdl_arr_6,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
input 	tdl_arr_4;
output 	tdl_arr_6;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr~6_combout ;
wire \tdl_arr[0]~q ;
wire \tdl_arr~5_combout ;
wire \tdl_arr[1]~q ;
wire \tdl_arr~4_combout ;
wire \tdl_arr[2]~q ;
wire \tdl_arr~3_combout ;
wire \tdl_arr[3]~q ;
wire \tdl_arr~2_combout ;
wire \tdl_arr[4]~q ;
wire \tdl_arr~1_combout ;
wire \tdl_arr[5]~q ;
wire \tdl_arr~0_combout ;


dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(tdl_arr_6),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~6 (
	.dataa(reset_n),
	.datab(tdl_arr_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~6_combout ),
	.cout());
defparam \tdl_arr~6 .lut_mask = 16'hEEEE;
defparam \tdl_arr~6 .sum_lutc_input = "datac";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(\tdl_arr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~5 (
	.dataa(reset_n),
	.datab(\tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~5_combout ),
	.cout());
defparam \tdl_arr~5 .lut_mask = 16'hEEEE;
defparam \tdl_arr~5 .sum_lutc_input = "datac";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~4 (
	.dataa(reset_n),
	.datab(\tdl_arr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~4_combout ),
	.cout());
defparam \tdl_arr~4 .lut_mask = 16'hEEEE;
defparam \tdl_arr~4 .sum_lutc_input = "datac";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~3 (
	.dataa(reset_n),
	.datab(\tdl_arr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~3_combout ),
	.cout());
defparam \tdl_arr~3 .lut_mask = 16'hEEEE;
defparam \tdl_arr~3 .sum_lutc_input = "datac";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~2 (
	.dataa(reset_n),
	.datab(\tdl_arr[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~2_combout ),
	.cout());
defparam \tdl_arr~2 .lut_mask = 16'hEEEE;
defparam \tdl_arr~2 .sum_lutc_input = "datac";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~1 (
	.dataa(reset_n),
	.datab(\tdl_arr[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~1_combout ),
	.cout());
defparam \tdl_arr~1 .lut_mask = 16'hEEEE;
defparam \tdl_arr~1 .sum_lutc_input = "datac";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

cycloneive_lcell_comb \tdl_arr~0 (
	.dataa(reset_n),
	.datab(\tdl_arr[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tdl_arr~0_combout ),
	.cout());
defparam \tdl_arr~0 .lut_mask = 16'hEEEE;
defparam \tdl_arr~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_twadgen (
	ram_block3a2,
	ram_block3a3,
	ram_block3a0,
	ram_block3a1,
	ram_block3a01,
	ram_block3a11,
	ram_block3a21,
	ram_block3a31,
	ram_block3a4,
	ram_block3a5,
	global_clock_enable,
	p_2,
	p_0,
	p_1,
	k_count_4,
	k_count_2,
	Mux1,
	k_count_6,
	k_count_3,
	k_count_5,
	Mux0,
	k_count_7,
	Mux01,
	Mux11,
	Mux12,
	Mux02,
	Mux03,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block3a2;
output 	ram_block3a3;
output 	ram_block3a0;
output 	ram_block3a1;
output 	ram_block3a01;
output 	ram_block3a11;
output 	ram_block3a21;
output 	ram_block3a31;
output 	ram_block3a4;
output 	ram_block3a5;
input 	global_clock_enable;
input 	p_2;
input 	p_0;
input 	p_1;
input 	k_count_4;
input 	k_count_2;
input 	Mux1;
input 	k_count_6;
input 	k_count_3;
input 	k_count_5;
input 	Mux0;
input 	k_count_7;
output 	Mux01;
input 	Mux11;
input 	Mux12;
input 	Mux02;
input 	Mux03;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~1 ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~3 ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~5 ;
wire \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ;
wire \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux7~0_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~1 ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~3 ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~5 ;
wire \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1_combout ;
wire \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \Mux6~0_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux4~0_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;

wire [143:0] \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus ;
wire [143:0] \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus ;

assign ram_block3a2 = \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus [0];

assign ram_block3a3 = \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus [0];

assign ram_block3a0 = \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus [0];

assign ram_block3a1 = \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus [0];

assign ram_block3a01 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus [0];

assign ram_block3a11 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus [0];

assign ram_block3a21 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus [0];

assign ram_block3a31 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus [0];

assign ram_block3a4 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus [0];

assign ram_block3a5 = \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus [0];

cycloneive_ram_block \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_block3a0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_0|shift_taps_amm:auto_generated|altsyncram_4b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .operation_mode = "dual_port";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_first_bit_number = 2;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_first_bit_number = 2;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a2 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_block3a1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_0|shift_taps_amm:auto_generated|altsyncram_4b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .operation_mode = "dual_port";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_first_bit_number = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_first_bit_number = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a3 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux1~1_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_0|shift_taps_amm:auto_generated|altsyncram_4b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .operation_mode = "dual_port";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_bit_number = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_bit_number = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a0 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux0~2_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_0|shift_taps_amm:auto_generated|altsyncram_4b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .operation_mode = "dual_port";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_bit_number = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_width = 3;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_width = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_address = 0;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_bit_number = 1;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_last_address = 5;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_width = 4;
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_0|auto_generated|altsyncram2|ram_block3a1 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux7~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_first_bit_number = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_first_bit_number = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a0 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux6~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_first_bit_number = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_first_bit_number = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a1 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux5~1_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_first_bit_number = 2;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_first_bit_number = 2;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a2 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux4~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_first_bit_number = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_first_bit_number = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a3 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux3~3_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_first_bit_number = 4;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_first_bit_number = 4;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a4 .ram_block_type = "auto";

cycloneive_ram_block \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux2~3_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ,\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5_PORTBDATAOUT_bus ));
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_core_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_input_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .clk0_output_clock_enable = "ena0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .data_interleave_offset_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .data_interleave_width_in_bits = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_twadgen:twid_factors|altshift_taps:twad_temp_rtl_1|shift_taps_dmm:auto_generated|altsyncram_8b81:altsyncram2|ALTSYNCRAM";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .mixed_port_feed_through_mode = "old";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .operation_mode = "dual_port";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_out_clock = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_first_bit_number = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_address_width = 3;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_out_clear = "none";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_out_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_data_width = 1;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_first_address = 0;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_first_bit_number = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_last_address = 5;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_logical_ram_depth = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_logical_ram_width = 6;
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .port_b_read_enable_clock = "clock0";
defparam \twad_temp_rtl_1|auto_generated|altsyncram2|ram_block3a5 .ram_block_type = "auto";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(p_2),
	.datab(p_0),
	.datac(gnd),
	.datad(p_1),
	.cin(gnd),
	.combout(Mux01),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hEEFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ),
	.cout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~1 ));
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0 .lut_mask = 16'h55AA;
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~1 ),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ),
	.cout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~3 ));
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2 .lut_mask = 16'h5A5F;
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .lut_mask = 16'h7777;
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ),
	.datab(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.datac(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datad(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2_combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2 .lut_mask = 16'hFFFB;
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[1]~3 ),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ),
	.cout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~5 ));
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4 .lut_mask = 16'h5AAF;
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\twad_temp_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3_combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3 .lut_mask = 16'hAAFF;
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[2]~5 ),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6 .lut_mask = 16'hF0F0;
defparam \twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.datab(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datac(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 16'hFEFF;
defparam \twad_temp_rtl_0|auto_generated|cntr1|cout_actual .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 (
	.dataa(\twad_temp_rtl_0|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\twad_temp_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cout());
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .lut_mask = 16'hAAFF;
defparam \twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\twad_temp_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \twad_temp_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(k_count_6),
	.datab(Mux1),
	.datac(Mux01),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hEFFE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(Mux11),
	.datab(Mux12),
	.datac(p_1),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hEFFE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(k_count_7),
	.datab(Mux0),
	.datac(Mux01),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hEFFE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(Mux02),
	.datab(Mux03),
	.datac(p_1),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hEFFE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(p_0),
	.datab(k_count_6),
	.datac(p_2),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hEFFF;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ),
	.cout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~1 ));
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0 .lut_mask = 16'h55AA;
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~1 ),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ),
	.cout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~3 ));
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2 .lut_mask = 16'h5A5F;
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cout());
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0 .lut_mask = 16'hDDDD;
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~2_combout ),
	.datab(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.datac(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datad(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2_combout ),
	.cout());
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2 .lut_mask = 16'hFFBF;
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[1]~3 ),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ),
	.cout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~5 ));
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4 .lut_mask = 16'h5AAF;
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~4_combout ),
	.datab(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.datac(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datad(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3_combout ),
	.cout());
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3 .lut_mask = 16'hFFBF;
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[2]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[2]~5 ),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.cout());
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6 .lut_mask = 16'hF0F0;
defparam \twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1 (
	.dataa(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[0]~0_combout ),
	.datab(\twad_temp_rtl_1|auto_generated|cntr1|add_sub4_result_int[3]~6_combout ),
	.datac(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datad(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cin(gnd),
	.combout(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1_combout ),
	.cout());
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1 .lut_mask = 16'hFFBF;
defparam \twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1 .sum_lutc_input = "datac";

dffeas \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\twad_temp_rtl_1|auto_generated|cntr1|trigger_mux_w[0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \twad_temp_rtl_1|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(p_0),
	.datab(k_count_7),
	.datac(p_2),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hEFFF;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(gnd),
	.datab(p_0),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'h3CFF;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\Mux5~0_combout ),
	.datab(k_count_6),
	.datac(k_count_4),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFAFC;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(\Mux5~0_combout ),
	.datab(k_count_7),
	.datac(k_count_5),
	.datad(p_1),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hFAFC;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~2 (
	.dataa(k_count_6),
	.datab(k_count_2),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hACFF;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~3 (
	.dataa(p_1),
	.datab(p_0),
	.datac(Mux12),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
defparam \Mux3~3 .lut_mask = 16'hFFB8;
defparam \Mux3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(k_count_7),
	.datab(k_count_3),
	.datac(p_1),
	.datad(p_2),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hACFF;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~3 (
	.dataa(p_1),
	.datab(p_0),
	.datac(Mux03),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFFB8;
defparam \Mux2~3 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_unbburst_ctrl (
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_1,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_19,
	q_b_191,
	q_b_192,
	q_b_193,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_18,
	q_b_181,
	q_b_182,
	q_b_183,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_17,
	q_b_171,
	q_b_172,
	q_b_173,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_16,
	q_b_161,
	q_b_162,
	q_b_163,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_154,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_144,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	lpp_c_i,
	ram_in_reg_2_3,
	ram_in_reg_1_3,
	ram_in_reg_3_3,
	ram_in_reg_5_3,
	ram_block3a0,
	ram_block3a1,
	ram_in_reg_2_0,
	ram_in_reg_1_0,
	ram_in_reg_3_0,
	ram_in_reg_5_0,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_3_1,
	ram_in_reg_5_1,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_3_2,
	ram_in_reg_5_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_1_31,
	ram_in_reg_1_01,
	ram_in_reg_1_11,
	ram_in_reg_1_21,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	ram_in_reg_0_3,
	ram_in_reg_0_0,
	ram_in_reg_0_1,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	ram_in_reg_9_3,
	ram_in_reg_9_0,
	ram_in_reg_9_1,
	ram_in_reg_9_2,
	ram_in_reg_9_7,
	ram_in_reg_9_4,
	ram_in_reg_9_5,
	ram_in_reg_9_6,
	ram_in_reg_8_3,
	ram_in_reg_8_0,
	ram_in_reg_8_1,
	ram_in_reg_8_2,
	ram_in_reg_8_7,
	ram_in_reg_8_4,
	ram_in_reg_8_5,
	ram_in_reg_8_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_5_31,
	ram_in_reg_5_01,
	ram_in_reg_5_11,
	ram_in_reg_5_21,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_3_31,
	ram_in_reg_3_01,
	ram_in_reg_3_11,
	ram_in_reg_3_21,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	global_clock_enable,
	a_ram_data_in_bus_12,
	wraddress_a_bus_0,
	wraddress_a_bus_1,
	wraddress_a_bus_18,
	wraddress_a_bus_3,
	wraddress_a_bus_20,
	wraddress_a_bus_5,
	wraddress_a_bus_14,
	wraddress_a_bus_15,
	rdaddress_a_bus_0,
	rdaddress_a_bus_1,
	rdaddress_a_bus_18,
	rdaddress_a_bus_3,
	rdaddress_a_bus_20,
	rdaddress_a_bus_5,
	rdaddress_a_bus_22,
	rdaddress_a_bus_7,
	a_ram_data_in_bus_72,
	wraddress_a_bus_24,
	wraddress_a_bus_25,
	wraddress_a_bus_10,
	wraddress_a_bus_27,
	wraddress_a_bus_12,
	wraddress_a_bus_29,
	rdaddress_a_bus_24,
	rdaddress_a_bus_25,
	rdaddress_a_bus_10,
	rdaddress_a_bus_27,
	rdaddress_a_bus_12,
	rdaddress_a_bus_29,
	rdaddress_a_bus_14,
	rdaddress_a_bus_31,
	a_ram_data_in_bus_52,
	wraddress_a_bus_17,
	wraddress_a_bus_19,
	wraddress_a_bus_21,
	rdaddress_a_bus_17,
	rdaddress_a_bus_19,
	rdaddress_a_bus_21,
	rdaddress_a_bus_23,
	a_ram_data_in_bus_32,
	wraddress_a_bus_9,
	wraddress_a_bus_11,
	wraddress_a_bus_13,
	rdaddress_a_bus_9,
	rdaddress_a_bus_11,
	rdaddress_a_bus_13,
	rdaddress_a_bus_15,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_62,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_71,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_70,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_30,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_79,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_69,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_78,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_68,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_17,
	a_ram_data_in_bus_77,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_67,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_76,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_66,
	a_ram_data_in_bus_46,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_75,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_65,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_14,
	a_ram_data_in_bus_74,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_64,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_73,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_23,
	wc_vec_3,
	data_in_r_2,
	sel_ram_in,
	ram_in_reg_0_11,
	wr_address_i_int_0,
	data_rdy_vec_2,
	wr_address_i_int_1,
	ram_in_reg_2_11,
	wr_address_i_int_2,
	wr_address_i_int_3,
	ram_in_reg_4_11,
	wr_address_i_int_4,
	wr_address_i_int_5,
	wr_address_i_int_6,
	wr_address_i_int_7,
	ram_in_reg_0_12,
	ram_in_reg_0_01,
	data_rdy_vec_0,
	ram_in_reg_1_32,
	ram_in_reg_1_02,
	ram_in_reg_2_12,
	ram_in_reg_2_01,
	ram_in_reg_3_32,
	ram_in_reg_3_02,
	ram_in_reg_4_12,
	ram_in_reg_4_01,
	ram_in_reg_5_32,
	ram_in_reg_5_02,
	ram_in_reg_6_01,
	ram_in_reg_6_11,
	ram_in_reg_7_01,
	ram_in_reg_7_31,
	ram_in_reg_0_02,
	ram_in_reg_2_02,
	ram_in_reg_4_02,
	ram_in_reg_0_03,
	ram_in_reg_1_03,
	ram_in_reg_2_03,
	ram_in_reg_3_03,
	ram_in_reg_4_03,
	ram_in_reg_5_03,
	ram_in_reg_7_21,
	ram_in_reg_1_12,
	ram_in_reg_3_12,
	ram_in_reg_5_12,
	ram_in_reg_1_22,
	ram_in_reg_3_22,
	ram_in_reg_5_22,
	data_in_i_2,
	data_in_r_1,
	data_in_i_1,
	data_in_r_0,
	data_in_i_0,
	data_in_r_9,
	data_in_i_9,
	data_in_r_8,
	data_in_i_8,
	data_in_r_7,
	data_in_i_7,
	data_in_r_6,
	data_in_i_6,
	data_in_r_5,
	data_in_i_5,
	data_in_r_4,
	data_in_i_4,
	data_in_r_3,
	data_in_i_3,
	ram_data_out0_17,
	ram_data_out1_17,
	ram_data_out2_17,
	ram_data_out3_17,
	ram_data_out0_15,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_16,
	ram_data_out1_16,
	ram_data_out2_16,
	ram_data_out3_16,
	ram_data_out0_18,
	ram_data_out1_18,
	ram_data_out2_18,
	ram_data_out3_18,
	ram_data_out0_14,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_13,
	ram_data_out1_13,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_12,
	ram_data_out1_12,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_11,
	ram_data_out1_11,
	ram_data_out2_10,
	ram_data_out3_10,
	ram_data_out0_10,
	ram_data_out1_10,
	ram_data_out0_19,
	ram_data_out1_19,
	ram_data_out2_19,
	ram_data_out3_19,
	ram_data_out0_5,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_6,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_7,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_4,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_3,
	ram_data_out1_3,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_2,
	ram_data_out1_2,
	ram_data_out2_1,
	ram_data_out3_1,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_0,
	ram_data_out3_0,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out2_9,
	ram_data_out3_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	q_b_12;
input 	q_b_121;
input 	q_b_122;
input 	q_b_123;
input 	q_b_2;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_11;
input 	q_b_111;
input 	q_b_112;
input 	q_b_113;
input 	q_b_1;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_10;
input 	q_b_101;
input 	q_b_102;
input 	q_b_103;
input 	q_b_0;
input 	q_b_01;
input 	q_b_02;
input 	q_b_03;
input 	q_b_19;
input 	q_b_191;
input 	q_b_192;
input 	q_b_193;
input 	q_b_9;
input 	q_b_91;
input 	q_b_92;
input 	q_b_93;
input 	q_b_18;
input 	q_b_181;
input 	q_b_182;
input 	q_b_183;
input 	q_b_8;
input 	q_b_81;
input 	q_b_82;
input 	q_b_83;
input 	q_b_17;
input 	q_b_171;
input 	q_b_172;
input 	q_b_173;
input 	q_b_7;
input 	q_b_71;
input 	q_b_72;
input 	q_b_73;
input 	q_b_16;
input 	q_b_161;
input 	q_b_162;
input 	q_b_163;
input 	q_b_6;
input 	q_b_61;
input 	q_b_62;
input 	q_b_63;
input 	q_b_151;
input 	q_b_152;
input 	q_b_153;
input 	q_b_154;
input 	q_b_5;
input 	q_b_51;
input 	q_b_52;
input 	q_b_53;
input 	q_b_141;
input 	q_b_142;
input 	q_b_143;
input 	q_b_144;
input 	q_b_4;
input 	q_b_41;
input 	q_b_42;
input 	q_b_43;
input 	q_b_131;
input 	q_b_132;
input 	q_b_133;
input 	q_b_134;
input 	q_b_3;
input 	q_b_31;
input 	q_b_32;
input 	q_b_33;
input 	lpp_c_i;
input 	ram_in_reg_2_3;
input 	ram_in_reg_1_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_5_3;
input 	ram_block3a0;
input 	ram_block3a1;
input 	ram_in_reg_2_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_6;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_0;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_6;
input 	ram_in_reg_9_3;
input 	ram_in_reg_9_0;
input 	ram_in_reg_9_1;
input 	ram_in_reg_9_2;
input 	ram_in_reg_9_7;
input 	ram_in_reg_9_4;
input 	ram_in_reg_9_5;
input 	ram_in_reg_9_6;
input 	ram_in_reg_8_3;
input 	ram_in_reg_8_0;
input 	ram_in_reg_8_1;
input 	ram_in_reg_8_2;
input 	ram_in_reg_8_7;
input 	ram_in_reg_8_4;
input 	ram_in_reg_8_5;
input 	ram_in_reg_8_6;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_6;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_6;
input 	ram_in_reg_5_31;
input 	ram_in_reg_5_01;
input 	ram_in_reg_5_11;
input 	ram_in_reg_5_21;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_6;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_6;
input 	ram_in_reg_3_31;
input 	ram_in_reg_3_01;
input 	ram_in_reg_3_11;
input 	ram_in_reg_3_21;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_6;
input 	global_clock_enable;
output 	a_ram_data_in_bus_12;
output 	wraddress_a_bus_0;
output 	wraddress_a_bus_1;
output 	wraddress_a_bus_18;
output 	wraddress_a_bus_3;
output 	wraddress_a_bus_20;
output 	wraddress_a_bus_5;
output 	wraddress_a_bus_14;
output 	wraddress_a_bus_15;
output 	rdaddress_a_bus_0;
output 	rdaddress_a_bus_1;
output 	rdaddress_a_bus_18;
output 	rdaddress_a_bus_3;
output 	rdaddress_a_bus_20;
output 	rdaddress_a_bus_5;
output 	rdaddress_a_bus_22;
output 	rdaddress_a_bus_7;
output 	a_ram_data_in_bus_72;
output 	wraddress_a_bus_24;
output 	wraddress_a_bus_25;
output 	wraddress_a_bus_10;
output 	wraddress_a_bus_27;
output 	wraddress_a_bus_12;
output 	wraddress_a_bus_29;
output 	rdaddress_a_bus_24;
output 	rdaddress_a_bus_25;
output 	rdaddress_a_bus_10;
output 	rdaddress_a_bus_27;
output 	rdaddress_a_bus_12;
output 	rdaddress_a_bus_29;
output 	rdaddress_a_bus_14;
output 	rdaddress_a_bus_31;
output 	a_ram_data_in_bus_52;
output 	wraddress_a_bus_17;
output 	wraddress_a_bus_19;
output 	wraddress_a_bus_21;
output 	rdaddress_a_bus_17;
output 	rdaddress_a_bus_19;
output 	rdaddress_a_bus_21;
output 	rdaddress_a_bus_23;
output 	a_ram_data_in_bus_32;
output 	wraddress_a_bus_9;
output 	wraddress_a_bus_11;
output 	wraddress_a_bus_13;
output 	rdaddress_a_bus_9;
output 	rdaddress_a_bus_11;
output 	rdaddress_a_bus_13;
output 	rdaddress_a_bus_15;
output 	a_ram_data_in_bus_2;
output 	a_ram_data_in_bus_62;
output 	a_ram_data_in_bus_42;
output 	a_ram_data_in_bus_22;
output 	a_ram_data_in_bus_11;
output 	a_ram_data_in_bus_71;
output 	a_ram_data_in_bus_51;
output 	a_ram_data_in_bus_31;
output 	a_ram_data_in_bus_1;
output 	a_ram_data_in_bus_61;
output 	a_ram_data_in_bus_41;
output 	a_ram_data_in_bus_21;
output 	a_ram_data_in_bus_10;
output 	a_ram_data_in_bus_70;
output 	a_ram_data_in_bus_50;
output 	a_ram_data_in_bus_30;
output 	a_ram_data_in_bus_0;
output 	a_ram_data_in_bus_60;
output 	a_ram_data_in_bus_40;
output 	a_ram_data_in_bus_20;
output 	a_ram_data_in_bus_19;
output 	a_ram_data_in_bus_79;
output 	a_ram_data_in_bus_59;
output 	a_ram_data_in_bus_39;
output 	a_ram_data_in_bus_9;
output 	a_ram_data_in_bus_69;
output 	a_ram_data_in_bus_49;
output 	a_ram_data_in_bus_29;
output 	a_ram_data_in_bus_18;
output 	a_ram_data_in_bus_78;
output 	a_ram_data_in_bus_58;
output 	a_ram_data_in_bus_38;
output 	a_ram_data_in_bus_8;
output 	a_ram_data_in_bus_68;
output 	a_ram_data_in_bus_48;
output 	a_ram_data_in_bus_28;
output 	a_ram_data_in_bus_17;
output 	a_ram_data_in_bus_77;
output 	a_ram_data_in_bus_57;
output 	a_ram_data_in_bus_37;
output 	a_ram_data_in_bus_7;
output 	a_ram_data_in_bus_67;
output 	a_ram_data_in_bus_47;
output 	a_ram_data_in_bus_27;
output 	a_ram_data_in_bus_16;
output 	a_ram_data_in_bus_76;
output 	a_ram_data_in_bus_56;
output 	a_ram_data_in_bus_36;
output 	a_ram_data_in_bus_6;
output 	a_ram_data_in_bus_66;
output 	a_ram_data_in_bus_46;
output 	a_ram_data_in_bus_26;
output 	a_ram_data_in_bus_15;
output 	a_ram_data_in_bus_75;
output 	a_ram_data_in_bus_55;
output 	a_ram_data_in_bus_35;
output 	a_ram_data_in_bus_5;
output 	a_ram_data_in_bus_65;
output 	a_ram_data_in_bus_45;
output 	a_ram_data_in_bus_25;
output 	a_ram_data_in_bus_14;
output 	a_ram_data_in_bus_74;
output 	a_ram_data_in_bus_54;
output 	a_ram_data_in_bus_34;
output 	a_ram_data_in_bus_4;
output 	a_ram_data_in_bus_64;
output 	a_ram_data_in_bus_44;
output 	a_ram_data_in_bus_24;
output 	a_ram_data_in_bus_13;
output 	a_ram_data_in_bus_73;
output 	a_ram_data_in_bus_53;
output 	a_ram_data_in_bus_33;
output 	a_ram_data_in_bus_3;
output 	a_ram_data_in_bus_63;
output 	a_ram_data_in_bus_43;
output 	a_ram_data_in_bus_23;
input 	wc_vec_3;
input 	data_in_r_2;
input 	sel_ram_in;
input 	ram_in_reg_0_11;
input 	wr_address_i_int_0;
input 	data_rdy_vec_2;
input 	wr_address_i_int_1;
input 	ram_in_reg_2_11;
input 	wr_address_i_int_2;
input 	wr_address_i_int_3;
input 	ram_in_reg_4_11;
input 	wr_address_i_int_4;
input 	wr_address_i_int_5;
input 	wr_address_i_int_6;
input 	wr_address_i_int_7;
input 	ram_in_reg_0_12;
input 	ram_in_reg_0_01;
input 	data_rdy_vec_0;
input 	ram_in_reg_1_32;
input 	ram_in_reg_1_02;
input 	ram_in_reg_2_12;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_32;
input 	ram_in_reg_3_02;
input 	ram_in_reg_4_12;
input 	ram_in_reg_4_01;
input 	ram_in_reg_5_32;
input 	ram_in_reg_5_02;
input 	ram_in_reg_6_01;
input 	ram_in_reg_6_11;
input 	ram_in_reg_7_01;
input 	ram_in_reg_7_31;
input 	ram_in_reg_0_02;
input 	ram_in_reg_2_02;
input 	ram_in_reg_4_02;
input 	ram_in_reg_0_03;
input 	ram_in_reg_1_03;
input 	ram_in_reg_2_03;
input 	ram_in_reg_3_03;
input 	ram_in_reg_4_03;
input 	ram_in_reg_5_03;
input 	ram_in_reg_7_21;
input 	ram_in_reg_1_12;
input 	ram_in_reg_3_12;
input 	ram_in_reg_5_12;
input 	ram_in_reg_1_22;
input 	ram_in_reg_3_22;
input 	ram_in_reg_5_22;
input 	data_in_i_2;
input 	data_in_r_1;
input 	data_in_i_1;
input 	data_in_r_0;
input 	data_in_i_0;
input 	data_in_r_9;
input 	data_in_i_9;
input 	data_in_r_8;
input 	data_in_i_8;
input 	data_in_r_7;
input 	data_in_i_7;
input 	data_in_r_6;
input 	data_in_i_6;
input 	data_in_r_5;
input 	data_in_i_5;
input 	data_in_r_4;
input 	data_in_i_4;
input 	data_in_r_3;
input 	data_in_i_3;
output 	ram_data_out0_17;
output 	ram_data_out1_17;
output 	ram_data_out2_17;
output 	ram_data_out3_17;
output 	ram_data_out0_15;
output 	ram_data_out1_15;
output 	ram_data_out2_15;
output 	ram_data_out3_15;
output 	ram_data_out0_16;
output 	ram_data_out1_16;
output 	ram_data_out2_16;
output 	ram_data_out3_16;
output 	ram_data_out0_18;
output 	ram_data_out1_18;
output 	ram_data_out2_18;
output 	ram_data_out3_18;
output 	ram_data_out0_14;
output 	ram_data_out1_14;
output 	ram_data_out2_14;
output 	ram_data_out3_14;
output 	ram_data_out2_13;
output 	ram_data_out3_13;
output 	ram_data_out0_13;
output 	ram_data_out1_13;
output 	ram_data_out2_12;
output 	ram_data_out3_12;
output 	ram_data_out0_12;
output 	ram_data_out1_12;
output 	ram_data_out2_11;
output 	ram_data_out3_11;
output 	ram_data_out0_11;
output 	ram_data_out1_11;
output 	ram_data_out2_10;
output 	ram_data_out3_10;
output 	ram_data_out0_10;
output 	ram_data_out1_10;
output 	ram_data_out0_19;
output 	ram_data_out1_19;
output 	ram_data_out2_19;
output 	ram_data_out3_19;
output 	ram_data_out0_5;
output 	ram_data_out1_5;
output 	ram_data_out2_5;
output 	ram_data_out3_5;
output 	ram_data_out0_6;
output 	ram_data_out1_6;
output 	ram_data_out2_6;
output 	ram_data_out3_6;
output 	ram_data_out0_7;
output 	ram_data_out1_7;
output 	ram_data_out2_7;
output 	ram_data_out3_7;
output 	ram_data_out0_8;
output 	ram_data_out1_8;
output 	ram_data_out2_8;
output 	ram_data_out3_8;
output 	ram_data_out0_4;
output 	ram_data_out1_4;
output 	ram_data_out2_4;
output 	ram_data_out3_4;
output 	ram_data_out2_3;
output 	ram_data_out3_3;
output 	ram_data_out0_3;
output 	ram_data_out1_3;
output 	ram_data_out2_2;
output 	ram_data_out3_2;
output 	ram_data_out0_2;
output 	ram_data_out1_2;
output 	ram_data_out2_1;
output 	ram_data_out3_1;
output 	ram_data_out0_1;
output 	ram_data_out1_1;
output 	ram_data_out2_0;
output 	ram_data_out3_0;
output 	ram_data_out0_0;
output 	ram_data_out1_0;
output 	ram_data_out0_9;
output 	ram_data_out1_9;
output 	ram_data_out2_9;
output 	ram_data_out3_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a_ram_data_in_bus~0_combout ;
wire \wraddress_a_bus~0_combout ;
wire \wraddress_a_bus~1_combout ;
wire \wraddress_a_bus~2_combout ;
wire \wraddress_a_bus~3_combout ;
wire \wraddress_a_bus~4_combout ;
wire \wraddress_a_bus~5_combout ;
wire \wraddress_a_bus~6_combout ;
wire \wraddress_a_bus~7_combout ;
wire \rdaddress_a_bus~0_combout ;
wire \rdaddress_a_bus~1_combout ;
wire \rdaddress_a_bus~2_combout ;
wire \rdaddress_a_bus~3_combout ;
wire \rdaddress_a_bus~4_combout ;
wire \rdaddress_a_bus~5_combout ;
wire \rdaddress_a_bus~6_combout ;
wire \rdaddress_a_bus~7_combout ;
wire \a_ram_data_in_bus~1_combout ;
wire \wraddress_a_bus~8_combout ;
wire \wraddress_a_bus~9_combout ;
wire \wraddress_a_bus~10_combout ;
wire \wraddress_a_bus~11_combout ;
wire \wraddress_a_bus~12_combout ;
wire \wraddress_a_bus~13_combout ;
wire \rdaddress_a_bus~8_combout ;
wire \rdaddress_a_bus~9_combout ;
wire \rdaddress_a_bus~10_combout ;
wire \rdaddress_a_bus~11_combout ;
wire \rdaddress_a_bus~12_combout ;
wire \rdaddress_a_bus~13_combout ;
wire \rdaddress_a_bus~14_combout ;
wire \rdaddress_a_bus~15_combout ;
wire \a_ram_data_in_bus~2_combout ;
wire \wraddress_a_bus~14_combout ;
wire \wraddress_a_bus~15_combout ;
wire \wraddress_a_bus~16_combout ;
wire \rdaddress_a_bus~16_combout ;
wire \rdaddress_a_bus~17_combout ;
wire \rdaddress_a_bus~18_combout ;
wire \rdaddress_a_bus~19_combout ;
wire \a_ram_data_in_bus~3_combout ;
wire \wraddress_a_bus~17_combout ;
wire \wraddress_a_bus~18_combout ;
wire \wraddress_a_bus~19_combout ;
wire \rdaddress_a_bus~20_combout ;
wire \rdaddress_a_bus~21_combout ;
wire \rdaddress_a_bus~22_combout ;
wire \rdaddress_a_bus~23_combout ;
wire \a_ram_data_in_bus~4_combout ;
wire \a_ram_data_in_bus~5_combout ;
wire \a_ram_data_in_bus~6_combout ;
wire \a_ram_data_in_bus~7_combout ;
wire \a_ram_data_in_bus~8_combout ;
wire \a_ram_data_in_bus~9_combout ;
wire \a_ram_data_in_bus~10_combout ;
wire \a_ram_data_in_bus~11_combout ;
wire \a_ram_data_in_bus~12_combout ;
wire \a_ram_data_in_bus~13_combout ;
wire \a_ram_data_in_bus~14_combout ;
wire \a_ram_data_in_bus~15_combout ;
wire \a_ram_data_in_bus~16_combout ;
wire \a_ram_data_in_bus~17_combout ;
wire \a_ram_data_in_bus~18_combout ;
wire \a_ram_data_in_bus~19_combout ;
wire \a_ram_data_in_bus~20_combout ;
wire \a_ram_data_in_bus~21_combout ;
wire \a_ram_data_in_bus~22_combout ;
wire \a_ram_data_in_bus~23_combout ;
wire \a_ram_data_in_bus~24_combout ;
wire \a_ram_data_in_bus~25_combout ;
wire \a_ram_data_in_bus~26_combout ;
wire \a_ram_data_in_bus~27_combout ;
wire \a_ram_data_in_bus~28_combout ;
wire \a_ram_data_in_bus~29_combout ;
wire \a_ram_data_in_bus~30_combout ;
wire \a_ram_data_in_bus~31_combout ;
wire \a_ram_data_in_bus~32_combout ;
wire \a_ram_data_in_bus~33_combout ;
wire \a_ram_data_in_bus~34_combout ;
wire \a_ram_data_in_bus~35_combout ;
wire \a_ram_data_in_bus~36_combout ;
wire \a_ram_data_in_bus~37_combout ;
wire \a_ram_data_in_bus~38_combout ;
wire \a_ram_data_in_bus~39_combout ;
wire \a_ram_data_in_bus~40_combout ;
wire \a_ram_data_in_bus~41_combout ;
wire \a_ram_data_in_bus~42_combout ;
wire \a_ram_data_in_bus~43_combout ;
wire \a_ram_data_in_bus~44_combout ;
wire \a_ram_data_in_bus~45_combout ;
wire \a_ram_data_in_bus~46_combout ;
wire \a_ram_data_in_bus~47_combout ;
wire \a_ram_data_in_bus~48_combout ;
wire \a_ram_data_in_bus~49_combout ;
wire \a_ram_data_in_bus~50_combout ;
wire \a_ram_data_in_bus~51_combout ;
wire \a_ram_data_in_bus~52_combout ;
wire \a_ram_data_in_bus~53_combout ;
wire \a_ram_data_in_bus~54_combout ;
wire \a_ram_data_in_bus~55_combout ;
wire \a_ram_data_in_bus~56_combout ;
wire \a_ram_data_in_bus~57_combout ;
wire \a_ram_data_in_bus~58_combout ;
wire \a_ram_data_in_bus~59_combout ;
wire \a_ram_data_in_bus~60_combout ;
wire \a_ram_data_in_bus~61_combout ;
wire \a_ram_data_in_bus~62_combout ;
wire \a_ram_data_in_bus~63_combout ;
wire \a_ram_data_in_bus~64_combout ;
wire \a_ram_data_in_bus~65_combout ;
wire \a_ram_data_in_bus~66_combout ;
wire \a_ram_data_in_bus~67_combout ;
wire \a_ram_data_in_bus~68_combout ;
wire \a_ram_data_in_bus~69_combout ;
wire \a_ram_data_in_bus~70_combout ;
wire \a_ram_data_in_bus~71_combout ;
wire \a_ram_data_in_bus~72_combout ;
wire \a_ram_data_in_bus~73_combout ;
wire \a_ram_data_in_bus~74_combout ;
wire \a_ram_data_in_bus~75_combout ;
wire \a_ram_data_in_bus~76_combout ;
wire \a_ram_data_in_bus~77_combout ;
wire \a_ram_data_in_bus~78_combout ;
wire \a_ram_data_in_bus~79_combout ;


dffeas \a_ram_data_in_bus[12] (
	.clk(clk),
	.d(\a_ram_data_in_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_12),
	.prn(vcc));
defparam \a_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[12] .power_up = "low";

dffeas \wraddress_a_bus[0] (
	.clk(clk),
	.d(\wraddress_a_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_0),
	.prn(vcc));
defparam \wraddress_a_bus[0] .is_wysiwyg = "true";
defparam \wraddress_a_bus[0] .power_up = "low";

dffeas \wraddress_a_bus[1] (
	.clk(clk),
	.d(\wraddress_a_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_1),
	.prn(vcc));
defparam \wraddress_a_bus[1] .is_wysiwyg = "true";
defparam \wraddress_a_bus[1] .power_up = "low";

dffeas \wraddress_a_bus[18] (
	.clk(clk),
	.d(\wraddress_a_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_18),
	.prn(vcc));
defparam \wraddress_a_bus[18] .is_wysiwyg = "true";
defparam \wraddress_a_bus[18] .power_up = "low";

dffeas \wraddress_a_bus[3] (
	.clk(clk),
	.d(\wraddress_a_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_3),
	.prn(vcc));
defparam \wraddress_a_bus[3] .is_wysiwyg = "true";
defparam \wraddress_a_bus[3] .power_up = "low";

dffeas \wraddress_a_bus[20] (
	.clk(clk),
	.d(\wraddress_a_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_20),
	.prn(vcc));
defparam \wraddress_a_bus[20] .is_wysiwyg = "true";
defparam \wraddress_a_bus[20] .power_up = "low";

dffeas \wraddress_a_bus[5] (
	.clk(clk),
	.d(\wraddress_a_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_5),
	.prn(vcc));
defparam \wraddress_a_bus[5] .is_wysiwyg = "true";
defparam \wraddress_a_bus[5] .power_up = "low";

dffeas \wraddress_a_bus[14] (
	.clk(clk),
	.d(\wraddress_a_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_14),
	.prn(vcc));
defparam \wraddress_a_bus[14] .is_wysiwyg = "true";
defparam \wraddress_a_bus[14] .power_up = "low";

dffeas \wraddress_a_bus[15] (
	.clk(clk),
	.d(\wraddress_a_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_15),
	.prn(vcc));
defparam \wraddress_a_bus[15] .is_wysiwyg = "true";
defparam \wraddress_a_bus[15] .power_up = "low";

dffeas \rdaddress_a_bus[0] (
	.clk(clk),
	.d(\rdaddress_a_bus~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_0),
	.prn(vcc));
defparam \rdaddress_a_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[0] .power_up = "low";

dffeas \rdaddress_a_bus[1] (
	.clk(clk),
	.d(\rdaddress_a_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_1),
	.prn(vcc));
defparam \rdaddress_a_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[1] .power_up = "low";

dffeas \rdaddress_a_bus[18] (
	.clk(clk),
	.d(\rdaddress_a_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_18),
	.prn(vcc));
defparam \rdaddress_a_bus[18] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[18] .power_up = "low";

dffeas \rdaddress_a_bus[3] (
	.clk(clk),
	.d(\rdaddress_a_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_3),
	.prn(vcc));
defparam \rdaddress_a_bus[3] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[3] .power_up = "low";

dffeas \rdaddress_a_bus[20] (
	.clk(clk),
	.d(\rdaddress_a_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_20),
	.prn(vcc));
defparam \rdaddress_a_bus[20] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[20] .power_up = "low";

dffeas \rdaddress_a_bus[5] (
	.clk(clk),
	.d(\rdaddress_a_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_5),
	.prn(vcc));
defparam \rdaddress_a_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[5] .power_up = "low";

dffeas \rdaddress_a_bus[22] (
	.clk(clk),
	.d(\rdaddress_a_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_22),
	.prn(vcc));
defparam \rdaddress_a_bus[22] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[22] .power_up = "low";

dffeas \rdaddress_a_bus[7] (
	.clk(clk),
	.d(\rdaddress_a_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_7),
	.prn(vcc));
defparam \rdaddress_a_bus[7] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[72] (
	.clk(clk),
	.d(\a_ram_data_in_bus~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_72),
	.prn(vcc));
defparam \a_ram_data_in_bus[72] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[72] .power_up = "low";

dffeas \wraddress_a_bus[24] (
	.clk(clk),
	.d(\wraddress_a_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_24),
	.prn(vcc));
defparam \wraddress_a_bus[24] .is_wysiwyg = "true";
defparam \wraddress_a_bus[24] .power_up = "low";

dffeas \wraddress_a_bus[25] (
	.clk(clk),
	.d(\wraddress_a_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_25),
	.prn(vcc));
defparam \wraddress_a_bus[25] .is_wysiwyg = "true";
defparam \wraddress_a_bus[25] .power_up = "low";

dffeas \wraddress_a_bus[10] (
	.clk(clk),
	.d(\wraddress_a_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_10),
	.prn(vcc));
defparam \wraddress_a_bus[10] .is_wysiwyg = "true";
defparam \wraddress_a_bus[10] .power_up = "low";

dffeas \wraddress_a_bus[27] (
	.clk(clk),
	.d(\wraddress_a_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_27),
	.prn(vcc));
defparam \wraddress_a_bus[27] .is_wysiwyg = "true";
defparam \wraddress_a_bus[27] .power_up = "low";

dffeas \wraddress_a_bus[12] (
	.clk(clk),
	.d(\wraddress_a_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_12),
	.prn(vcc));
defparam \wraddress_a_bus[12] .is_wysiwyg = "true";
defparam \wraddress_a_bus[12] .power_up = "low";

dffeas \wraddress_a_bus[29] (
	.clk(clk),
	.d(\wraddress_a_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_29),
	.prn(vcc));
defparam \wraddress_a_bus[29] .is_wysiwyg = "true";
defparam \wraddress_a_bus[29] .power_up = "low";

dffeas \rdaddress_a_bus[24] (
	.clk(clk),
	.d(\rdaddress_a_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_24),
	.prn(vcc));
defparam \rdaddress_a_bus[24] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[24] .power_up = "low";

dffeas \rdaddress_a_bus[25] (
	.clk(clk),
	.d(\rdaddress_a_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_25),
	.prn(vcc));
defparam \rdaddress_a_bus[25] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[25] .power_up = "low";

dffeas \rdaddress_a_bus[10] (
	.clk(clk),
	.d(\rdaddress_a_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_10),
	.prn(vcc));
defparam \rdaddress_a_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[10] .power_up = "low";

dffeas \rdaddress_a_bus[27] (
	.clk(clk),
	.d(\rdaddress_a_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_27),
	.prn(vcc));
defparam \rdaddress_a_bus[27] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[27] .power_up = "low";

dffeas \rdaddress_a_bus[12] (
	.clk(clk),
	.d(\rdaddress_a_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_12),
	.prn(vcc));
defparam \rdaddress_a_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[12] .power_up = "low";

dffeas \rdaddress_a_bus[29] (
	.clk(clk),
	.d(\rdaddress_a_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_29),
	.prn(vcc));
defparam \rdaddress_a_bus[29] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[29] .power_up = "low";

dffeas \rdaddress_a_bus[14] (
	.clk(clk),
	.d(\rdaddress_a_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_14),
	.prn(vcc));
defparam \rdaddress_a_bus[14] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[14] .power_up = "low";

dffeas \rdaddress_a_bus[31] (
	.clk(clk),
	.d(\rdaddress_a_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_31),
	.prn(vcc));
defparam \rdaddress_a_bus[31] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[31] .power_up = "low";

dffeas \a_ram_data_in_bus[52] (
	.clk(clk),
	.d(\a_ram_data_in_bus~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_52),
	.prn(vcc));
defparam \a_ram_data_in_bus[52] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[52] .power_up = "low";

dffeas \wraddress_a_bus[17] (
	.clk(clk),
	.d(\wraddress_a_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_17),
	.prn(vcc));
defparam \wraddress_a_bus[17] .is_wysiwyg = "true";
defparam \wraddress_a_bus[17] .power_up = "low";

dffeas \wraddress_a_bus[19] (
	.clk(clk),
	.d(\wraddress_a_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_19),
	.prn(vcc));
defparam \wraddress_a_bus[19] .is_wysiwyg = "true";
defparam \wraddress_a_bus[19] .power_up = "low";

dffeas \wraddress_a_bus[21] (
	.clk(clk),
	.d(\wraddress_a_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_21),
	.prn(vcc));
defparam \wraddress_a_bus[21] .is_wysiwyg = "true";
defparam \wraddress_a_bus[21] .power_up = "low";

dffeas \rdaddress_a_bus[17] (
	.clk(clk),
	.d(\rdaddress_a_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_17),
	.prn(vcc));
defparam \rdaddress_a_bus[17] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[17] .power_up = "low";

dffeas \rdaddress_a_bus[19] (
	.clk(clk),
	.d(\rdaddress_a_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_19),
	.prn(vcc));
defparam \rdaddress_a_bus[19] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[19] .power_up = "low";

dffeas \rdaddress_a_bus[21] (
	.clk(clk),
	.d(\rdaddress_a_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_21),
	.prn(vcc));
defparam \rdaddress_a_bus[21] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[21] .power_up = "low";

dffeas \rdaddress_a_bus[23] (
	.clk(clk),
	.d(\rdaddress_a_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_23),
	.prn(vcc));
defparam \rdaddress_a_bus[23] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[23] .power_up = "low";

dffeas \a_ram_data_in_bus[32] (
	.clk(clk),
	.d(\a_ram_data_in_bus~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_32),
	.prn(vcc));
defparam \a_ram_data_in_bus[32] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[32] .power_up = "low";

dffeas \wraddress_a_bus[9] (
	.clk(clk),
	.d(\wraddress_a_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_9),
	.prn(vcc));
defparam \wraddress_a_bus[9] .is_wysiwyg = "true";
defparam \wraddress_a_bus[9] .power_up = "low";

dffeas \wraddress_a_bus[11] (
	.clk(clk),
	.d(\wraddress_a_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_11),
	.prn(vcc));
defparam \wraddress_a_bus[11] .is_wysiwyg = "true";
defparam \wraddress_a_bus[11] .power_up = "low";

dffeas \wraddress_a_bus[13] (
	.clk(clk),
	.d(\wraddress_a_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(wraddress_a_bus_13),
	.prn(vcc));
defparam \wraddress_a_bus[13] .is_wysiwyg = "true";
defparam \wraddress_a_bus[13] .power_up = "low";

dffeas \rdaddress_a_bus[9] (
	.clk(clk),
	.d(\rdaddress_a_bus~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_9),
	.prn(vcc));
defparam \rdaddress_a_bus[9] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[9] .power_up = "low";

dffeas \rdaddress_a_bus[11] (
	.clk(clk),
	.d(\rdaddress_a_bus~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_11),
	.prn(vcc));
defparam \rdaddress_a_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[11] .power_up = "low";

dffeas \rdaddress_a_bus[13] (
	.clk(clk),
	.d(\rdaddress_a_bus~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_13),
	.prn(vcc));
defparam \rdaddress_a_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[13] .power_up = "low";

dffeas \rdaddress_a_bus[15] (
	.clk(clk),
	.d(\rdaddress_a_bus~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(rdaddress_a_bus_15),
	.prn(vcc));
defparam \rdaddress_a_bus[15] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[15] .power_up = "low";

dffeas \a_ram_data_in_bus[2] (
	.clk(clk),
	.d(\a_ram_data_in_bus~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_2),
	.prn(vcc));
defparam \a_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[2] .power_up = "low";

dffeas \a_ram_data_in_bus[62] (
	.clk(clk),
	.d(\a_ram_data_in_bus~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_62),
	.prn(vcc));
defparam \a_ram_data_in_bus[62] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[62] .power_up = "low";

dffeas \a_ram_data_in_bus[42] (
	.clk(clk),
	.d(\a_ram_data_in_bus~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_42),
	.prn(vcc));
defparam \a_ram_data_in_bus[42] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[42] .power_up = "low";

dffeas \a_ram_data_in_bus[22] (
	.clk(clk),
	.d(\a_ram_data_in_bus~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_22),
	.prn(vcc));
defparam \a_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[22] .power_up = "low";

dffeas \a_ram_data_in_bus[11] (
	.clk(clk),
	.d(\a_ram_data_in_bus~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_11),
	.prn(vcc));
defparam \a_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[11] .power_up = "low";

dffeas \a_ram_data_in_bus[71] (
	.clk(clk),
	.d(\a_ram_data_in_bus~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_71),
	.prn(vcc));
defparam \a_ram_data_in_bus[71] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[71] .power_up = "low";

dffeas \a_ram_data_in_bus[51] (
	.clk(clk),
	.d(\a_ram_data_in_bus~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_51),
	.prn(vcc));
defparam \a_ram_data_in_bus[51] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[51] .power_up = "low";

dffeas \a_ram_data_in_bus[31] (
	.clk(clk),
	.d(\a_ram_data_in_bus~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_31),
	.prn(vcc));
defparam \a_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[31] .power_up = "low";

dffeas \a_ram_data_in_bus[1] (
	.clk(clk),
	.d(\a_ram_data_in_bus~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_1),
	.prn(vcc));
defparam \a_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[1] .power_up = "low";

dffeas \a_ram_data_in_bus[61] (
	.clk(clk),
	.d(\a_ram_data_in_bus~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_61),
	.prn(vcc));
defparam \a_ram_data_in_bus[61] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[61] .power_up = "low";

dffeas \a_ram_data_in_bus[41] (
	.clk(clk),
	.d(\a_ram_data_in_bus~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_41),
	.prn(vcc));
defparam \a_ram_data_in_bus[41] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[41] .power_up = "low";

dffeas \a_ram_data_in_bus[21] (
	.clk(clk),
	.d(\a_ram_data_in_bus~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_21),
	.prn(vcc));
defparam \a_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[21] .power_up = "low";

dffeas \a_ram_data_in_bus[10] (
	.clk(clk),
	.d(\a_ram_data_in_bus~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_10),
	.prn(vcc));
defparam \a_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[10] .power_up = "low";

dffeas \a_ram_data_in_bus[70] (
	.clk(clk),
	.d(\a_ram_data_in_bus~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_70),
	.prn(vcc));
defparam \a_ram_data_in_bus[70] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[70] .power_up = "low";

dffeas \a_ram_data_in_bus[50] (
	.clk(clk),
	.d(\a_ram_data_in_bus~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_50),
	.prn(vcc));
defparam \a_ram_data_in_bus[50] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[50] .power_up = "low";

dffeas \a_ram_data_in_bus[30] (
	.clk(clk),
	.d(\a_ram_data_in_bus~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_30),
	.prn(vcc));
defparam \a_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[30] .power_up = "low";

dffeas \a_ram_data_in_bus[0] (
	.clk(clk),
	.d(\a_ram_data_in_bus~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_0),
	.prn(vcc));
defparam \a_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[0] .power_up = "low";

dffeas \a_ram_data_in_bus[60] (
	.clk(clk),
	.d(\a_ram_data_in_bus~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_60),
	.prn(vcc));
defparam \a_ram_data_in_bus[60] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[60] .power_up = "low";

dffeas \a_ram_data_in_bus[40] (
	.clk(clk),
	.d(\a_ram_data_in_bus~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_40),
	.prn(vcc));
defparam \a_ram_data_in_bus[40] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[40] .power_up = "low";

dffeas \a_ram_data_in_bus[20] (
	.clk(clk),
	.d(\a_ram_data_in_bus~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_20),
	.prn(vcc));
defparam \a_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[20] .power_up = "low";

dffeas \a_ram_data_in_bus[19] (
	.clk(clk),
	.d(\a_ram_data_in_bus~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_19),
	.prn(vcc));
defparam \a_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[19] .power_up = "low";

dffeas \a_ram_data_in_bus[79] (
	.clk(clk),
	.d(\a_ram_data_in_bus~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_79),
	.prn(vcc));
defparam \a_ram_data_in_bus[79] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[79] .power_up = "low";

dffeas \a_ram_data_in_bus[59] (
	.clk(clk),
	.d(\a_ram_data_in_bus~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_59),
	.prn(vcc));
defparam \a_ram_data_in_bus[59] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[59] .power_up = "low";

dffeas \a_ram_data_in_bus[39] (
	.clk(clk),
	.d(\a_ram_data_in_bus~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_39),
	.prn(vcc));
defparam \a_ram_data_in_bus[39] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[39] .power_up = "low";

dffeas \a_ram_data_in_bus[9] (
	.clk(clk),
	.d(\a_ram_data_in_bus~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_9),
	.prn(vcc));
defparam \a_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[9] .power_up = "low";

dffeas \a_ram_data_in_bus[69] (
	.clk(clk),
	.d(\a_ram_data_in_bus~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_69),
	.prn(vcc));
defparam \a_ram_data_in_bus[69] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[69] .power_up = "low";

dffeas \a_ram_data_in_bus[49] (
	.clk(clk),
	.d(\a_ram_data_in_bus~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_49),
	.prn(vcc));
defparam \a_ram_data_in_bus[49] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[49] .power_up = "low";

dffeas \a_ram_data_in_bus[29] (
	.clk(clk),
	.d(\a_ram_data_in_bus~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_29),
	.prn(vcc));
defparam \a_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[29] .power_up = "low";

dffeas \a_ram_data_in_bus[18] (
	.clk(clk),
	.d(\a_ram_data_in_bus~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_18),
	.prn(vcc));
defparam \a_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[18] .power_up = "low";

dffeas \a_ram_data_in_bus[78] (
	.clk(clk),
	.d(\a_ram_data_in_bus~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_78),
	.prn(vcc));
defparam \a_ram_data_in_bus[78] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[78] .power_up = "low";

dffeas \a_ram_data_in_bus[58] (
	.clk(clk),
	.d(\a_ram_data_in_bus~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_58),
	.prn(vcc));
defparam \a_ram_data_in_bus[58] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[58] .power_up = "low";

dffeas \a_ram_data_in_bus[38] (
	.clk(clk),
	.d(\a_ram_data_in_bus~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_38),
	.prn(vcc));
defparam \a_ram_data_in_bus[38] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[38] .power_up = "low";

dffeas \a_ram_data_in_bus[8] (
	.clk(clk),
	.d(\a_ram_data_in_bus~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_8),
	.prn(vcc));
defparam \a_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[8] .power_up = "low";

dffeas \a_ram_data_in_bus[68] (
	.clk(clk),
	.d(\a_ram_data_in_bus~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_68),
	.prn(vcc));
defparam \a_ram_data_in_bus[68] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[68] .power_up = "low";

dffeas \a_ram_data_in_bus[48] (
	.clk(clk),
	.d(\a_ram_data_in_bus~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_48),
	.prn(vcc));
defparam \a_ram_data_in_bus[48] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[48] .power_up = "low";

dffeas \a_ram_data_in_bus[28] (
	.clk(clk),
	.d(\a_ram_data_in_bus~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_28),
	.prn(vcc));
defparam \a_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[28] .power_up = "low";

dffeas \a_ram_data_in_bus[17] (
	.clk(clk),
	.d(\a_ram_data_in_bus~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_17),
	.prn(vcc));
defparam \a_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[17] .power_up = "low";

dffeas \a_ram_data_in_bus[77] (
	.clk(clk),
	.d(\a_ram_data_in_bus~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_77),
	.prn(vcc));
defparam \a_ram_data_in_bus[77] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[77] .power_up = "low";

dffeas \a_ram_data_in_bus[57] (
	.clk(clk),
	.d(\a_ram_data_in_bus~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_57),
	.prn(vcc));
defparam \a_ram_data_in_bus[57] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[57] .power_up = "low";

dffeas \a_ram_data_in_bus[37] (
	.clk(clk),
	.d(\a_ram_data_in_bus~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_37),
	.prn(vcc));
defparam \a_ram_data_in_bus[37] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[37] .power_up = "low";

dffeas \a_ram_data_in_bus[7] (
	.clk(clk),
	.d(\a_ram_data_in_bus~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_7),
	.prn(vcc));
defparam \a_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[67] (
	.clk(clk),
	.d(\a_ram_data_in_bus~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_67),
	.prn(vcc));
defparam \a_ram_data_in_bus[67] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[67] .power_up = "low";

dffeas \a_ram_data_in_bus[47] (
	.clk(clk),
	.d(\a_ram_data_in_bus~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_47),
	.prn(vcc));
defparam \a_ram_data_in_bus[47] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[47] .power_up = "low";

dffeas \a_ram_data_in_bus[27] (
	.clk(clk),
	.d(\a_ram_data_in_bus~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_27),
	.prn(vcc));
defparam \a_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[27] .power_up = "low";

dffeas \a_ram_data_in_bus[16] (
	.clk(clk),
	.d(\a_ram_data_in_bus~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_16),
	.prn(vcc));
defparam \a_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[16] .power_up = "low";

dffeas \a_ram_data_in_bus[76] (
	.clk(clk),
	.d(\a_ram_data_in_bus~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_76),
	.prn(vcc));
defparam \a_ram_data_in_bus[76] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[76] .power_up = "low";

dffeas \a_ram_data_in_bus[56] (
	.clk(clk),
	.d(\a_ram_data_in_bus~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_56),
	.prn(vcc));
defparam \a_ram_data_in_bus[56] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[56] .power_up = "low";

dffeas \a_ram_data_in_bus[36] (
	.clk(clk),
	.d(\a_ram_data_in_bus~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_36),
	.prn(vcc));
defparam \a_ram_data_in_bus[36] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[36] .power_up = "low";

dffeas \a_ram_data_in_bus[6] (
	.clk(clk),
	.d(\a_ram_data_in_bus~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_6),
	.prn(vcc));
defparam \a_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[6] .power_up = "low";

dffeas \a_ram_data_in_bus[66] (
	.clk(clk),
	.d(\a_ram_data_in_bus~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_66),
	.prn(vcc));
defparam \a_ram_data_in_bus[66] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[66] .power_up = "low";

dffeas \a_ram_data_in_bus[46] (
	.clk(clk),
	.d(\a_ram_data_in_bus~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_46),
	.prn(vcc));
defparam \a_ram_data_in_bus[46] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[46] .power_up = "low";

dffeas \a_ram_data_in_bus[26] (
	.clk(clk),
	.d(\a_ram_data_in_bus~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_26),
	.prn(vcc));
defparam \a_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[26] .power_up = "low";

dffeas \a_ram_data_in_bus[15] (
	.clk(clk),
	.d(\a_ram_data_in_bus~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_15),
	.prn(vcc));
defparam \a_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[15] .power_up = "low";

dffeas \a_ram_data_in_bus[75] (
	.clk(clk),
	.d(\a_ram_data_in_bus~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_75),
	.prn(vcc));
defparam \a_ram_data_in_bus[75] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[75] .power_up = "low";

dffeas \a_ram_data_in_bus[55] (
	.clk(clk),
	.d(\a_ram_data_in_bus~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_55),
	.prn(vcc));
defparam \a_ram_data_in_bus[55] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[55] .power_up = "low";

dffeas \a_ram_data_in_bus[35] (
	.clk(clk),
	.d(\a_ram_data_in_bus~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_35),
	.prn(vcc));
defparam \a_ram_data_in_bus[35] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[35] .power_up = "low";

dffeas \a_ram_data_in_bus[5] (
	.clk(clk),
	.d(\a_ram_data_in_bus~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_5),
	.prn(vcc));
defparam \a_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[65] (
	.clk(clk),
	.d(\a_ram_data_in_bus~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_65),
	.prn(vcc));
defparam \a_ram_data_in_bus[65] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[65] .power_up = "low";

dffeas \a_ram_data_in_bus[45] (
	.clk(clk),
	.d(\a_ram_data_in_bus~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_45),
	.prn(vcc));
defparam \a_ram_data_in_bus[45] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[45] .power_up = "low";

dffeas \a_ram_data_in_bus[25] (
	.clk(clk),
	.d(\a_ram_data_in_bus~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_25),
	.prn(vcc));
defparam \a_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[25] .power_up = "low";

dffeas \a_ram_data_in_bus[14] (
	.clk(clk),
	.d(\a_ram_data_in_bus~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_14),
	.prn(vcc));
defparam \a_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[14] .power_up = "low";

dffeas \a_ram_data_in_bus[74] (
	.clk(clk),
	.d(\a_ram_data_in_bus~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_74),
	.prn(vcc));
defparam \a_ram_data_in_bus[74] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[74] .power_up = "low";

dffeas \a_ram_data_in_bus[54] (
	.clk(clk),
	.d(\a_ram_data_in_bus~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_54),
	.prn(vcc));
defparam \a_ram_data_in_bus[54] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[54] .power_up = "low";

dffeas \a_ram_data_in_bus[34] (
	.clk(clk),
	.d(\a_ram_data_in_bus~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_34),
	.prn(vcc));
defparam \a_ram_data_in_bus[34] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[34] .power_up = "low";

dffeas \a_ram_data_in_bus[4] (
	.clk(clk),
	.d(\a_ram_data_in_bus~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_4),
	.prn(vcc));
defparam \a_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[4] .power_up = "low";

dffeas \a_ram_data_in_bus[64] (
	.clk(clk),
	.d(\a_ram_data_in_bus~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_64),
	.prn(vcc));
defparam \a_ram_data_in_bus[64] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[64] .power_up = "low";

dffeas \a_ram_data_in_bus[44] (
	.clk(clk),
	.d(\a_ram_data_in_bus~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_44),
	.prn(vcc));
defparam \a_ram_data_in_bus[44] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[44] .power_up = "low";

dffeas \a_ram_data_in_bus[24] (
	.clk(clk),
	.d(\a_ram_data_in_bus~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_24),
	.prn(vcc));
defparam \a_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[24] .power_up = "low";

dffeas \a_ram_data_in_bus[13] (
	.clk(clk),
	.d(\a_ram_data_in_bus~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_13),
	.prn(vcc));
defparam \a_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[73] (
	.clk(clk),
	.d(\a_ram_data_in_bus~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_73),
	.prn(vcc));
defparam \a_ram_data_in_bus[73] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[73] .power_up = "low";

dffeas \a_ram_data_in_bus[53] (
	.clk(clk),
	.d(\a_ram_data_in_bus~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_53),
	.prn(vcc));
defparam \a_ram_data_in_bus[53] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[53] .power_up = "low";

dffeas \a_ram_data_in_bus[33] (
	.clk(clk),
	.d(\a_ram_data_in_bus~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_33),
	.prn(vcc));
defparam \a_ram_data_in_bus[33] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[33] .power_up = "low";

dffeas \a_ram_data_in_bus[3] (
	.clk(clk),
	.d(\a_ram_data_in_bus~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_3),
	.prn(vcc));
defparam \a_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[3] .power_up = "low";

dffeas \a_ram_data_in_bus[63] (
	.clk(clk),
	.d(\a_ram_data_in_bus~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_63),
	.prn(vcc));
defparam \a_ram_data_in_bus[63] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[63] .power_up = "low";

dffeas \a_ram_data_in_bus[43] (
	.clk(clk),
	.d(\a_ram_data_in_bus~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_43),
	.prn(vcc));
defparam \a_ram_data_in_bus[43] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[43] .power_up = "low";

dffeas \a_ram_data_in_bus[23] (
	.clk(clk),
	.d(\a_ram_data_in_bus~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(a_ram_data_in_bus_23),
	.prn(vcc));
defparam \a_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[23] .power_up = "low";

dffeas \ram_data_out0[17] (
	.clk(clk),
	.d(q_b_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_17),
	.prn(vcc));
defparam \ram_data_out0[17] .is_wysiwyg = "true";
defparam \ram_data_out0[17] .power_up = "low";

dffeas \ram_data_out1[17] (
	.clk(clk),
	.d(q_b_172),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_17),
	.prn(vcc));
defparam \ram_data_out1[17] .is_wysiwyg = "true";
defparam \ram_data_out1[17] .power_up = "low";

dffeas \ram_data_out2[17] (
	.clk(clk),
	.d(q_b_173),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_17),
	.prn(vcc));
defparam \ram_data_out2[17] .is_wysiwyg = "true";
defparam \ram_data_out2[17] .power_up = "low";

dffeas \ram_data_out3[17] (
	.clk(clk),
	.d(q_b_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_17),
	.prn(vcc));
defparam \ram_data_out3[17] .is_wysiwyg = "true";
defparam \ram_data_out3[17] .power_up = "low";

dffeas \ram_data_out0[15] (
	.clk(clk),
	.d(q_b_152),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_15),
	.prn(vcc));
defparam \ram_data_out0[15] .is_wysiwyg = "true";
defparam \ram_data_out0[15] .power_up = "low";

dffeas \ram_data_out1[15] (
	.clk(clk),
	.d(q_b_153),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_15),
	.prn(vcc));
defparam \ram_data_out1[15] .is_wysiwyg = "true";
defparam \ram_data_out1[15] .power_up = "low";

dffeas \ram_data_out2[15] (
	.clk(clk),
	.d(q_b_154),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_15),
	.prn(vcc));
defparam \ram_data_out2[15] .is_wysiwyg = "true";
defparam \ram_data_out2[15] .power_up = "low";

dffeas \ram_data_out3[15] (
	.clk(clk),
	.d(q_b_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_15),
	.prn(vcc));
defparam \ram_data_out3[15] .is_wysiwyg = "true";
defparam \ram_data_out3[15] .power_up = "low";

dffeas \ram_data_out0[16] (
	.clk(clk),
	.d(q_b_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_16),
	.prn(vcc));
defparam \ram_data_out0[16] .is_wysiwyg = "true";
defparam \ram_data_out0[16] .power_up = "low";

dffeas \ram_data_out1[16] (
	.clk(clk),
	.d(q_b_162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_16),
	.prn(vcc));
defparam \ram_data_out1[16] .is_wysiwyg = "true";
defparam \ram_data_out1[16] .power_up = "low";

dffeas \ram_data_out2[16] (
	.clk(clk),
	.d(q_b_163),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_16),
	.prn(vcc));
defparam \ram_data_out2[16] .is_wysiwyg = "true";
defparam \ram_data_out2[16] .power_up = "low";

dffeas \ram_data_out3[16] (
	.clk(clk),
	.d(q_b_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_16),
	.prn(vcc));
defparam \ram_data_out3[16] .is_wysiwyg = "true";
defparam \ram_data_out3[16] .power_up = "low";

dffeas \ram_data_out0[18] (
	.clk(clk),
	.d(q_b_181),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_18),
	.prn(vcc));
defparam \ram_data_out0[18] .is_wysiwyg = "true";
defparam \ram_data_out0[18] .power_up = "low";

dffeas \ram_data_out1[18] (
	.clk(clk),
	.d(q_b_182),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_18),
	.prn(vcc));
defparam \ram_data_out1[18] .is_wysiwyg = "true";
defparam \ram_data_out1[18] .power_up = "low";

dffeas \ram_data_out2[18] (
	.clk(clk),
	.d(q_b_183),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_18),
	.prn(vcc));
defparam \ram_data_out2[18] .is_wysiwyg = "true";
defparam \ram_data_out2[18] .power_up = "low";

dffeas \ram_data_out3[18] (
	.clk(clk),
	.d(q_b_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_18),
	.prn(vcc));
defparam \ram_data_out3[18] .is_wysiwyg = "true";
defparam \ram_data_out3[18] .power_up = "low";

dffeas \ram_data_out0[14] (
	.clk(clk),
	.d(q_b_142),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_14),
	.prn(vcc));
defparam \ram_data_out0[14] .is_wysiwyg = "true";
defparam \ram_data_out0[14] .power_up = "low";

dffeas \ram_data_out1[14] (
	.clk(clk),
	.d(q_b_143),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_14),
	.prn(vcc));
defparam \ram_data_out1[14] .is_wysiwyg = "true";
defparam \ram_data_out1[14] .power_up = "low";

dffeas \ram_data_out2[14] (
	.clk(clk),
	.d(q_b_144),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_14),
	.prn(vcc));
defparam \ram_data_out2[14] .is_wysiwyg = "true";
defparam \ram_data_out2[14] .power_up = "low";

dffeas \ram_data_out3[14] (
	.clk(clk),
	.d(q_b_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_14),
	.prn(vcc));
defparam \ram_data_out3[14] .is_wysiwyg = "true";
defparam \ram_data_out3[14] .power_up = "low";

dffeas \ram_data_out2[13] (
	.clk(clk),
	.d(q_b_134),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_13),
	.prn(vcc));
defparam \ram_data_out2[13] .is_wysiwyg = "true";
defparam \ram_data_out2[13] .power_up = "low";

dffeas \ram_data_out3[13] (
	.clk(clk),
	.d(q_b_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_13),
	.prn(vcc));
defparam \ram_data_out3[13] .is_wysiwyg = "true";
defparam \ram_data_out3[13] .power_up = "low";

dffeas \ram_data_out0[13] (
	.clk(clk),
	.d(q_b_132),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_13),
	.prn(vcc));
defparam \ram_data_out0[13] .is_wysiwyg = "true";
defparam \ram_data_out0[13] .power_up = "low";

dffeas \ram_data_out1[13] (
	.clk(clk),
	.d(q_b_133),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_13),
	.prn(vcc));
defparam \ram_data_out1[13] .is_wysiwyg = "true";
defparam \ram_data_out1[13] .power_up = "low";

dffeas \ram_data_out2[12] (
	.clk(clk),
	.d(q_b_123),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_12),
	.prn(vcc));
defparam \ram_data_out2[12] .is_wysiwyg = "true";
defparam \ram_data_out2[12] .power_up = "low";

dffeas \ram_data_out3[12] (
	.clk(clk),
	.d(q_b_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_12),
	.prn(vcc));
defparam \ram_data_out3[12] .is_wysiwyg = "true";
defparam \ram_data_out3[12] .power_up = "low";

dffeas \ram_data_out0[12] (
	.clk(clk),
	.d(q_b_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_12),
	.prn(vcc));
defparam \ram_data_out0[12] .is_wysiwyg = "true";
defparam \ram_data_out0[12] .power_up = "low";

dffeas \ram_data_out1[12] (
	.clk(clk),
	.d(q_b_122),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_12),
	.prn(vcc));
defparam \ram_data_out1[12] .is_wysiwyg = "true";
defparam \ram_data_out1[12] .power_up = "low";

dffeas \ram_data_out2[11] (
	.clk(clk),
	.d(q_b_113),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_11),
	.prn(vcc));
defparam \ram_data_out2[11] .is_wysiwyg = "true";
defparam \ram_data_out2[11] .power_up = "low";

dffeas \ram_data_out3[11] (
	.clk(clk),
	.d(q_b_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_11),
	.prn(vcc));
defparam \ram_data_out3[11] .is_wysiwyg = "true";
defparam \ram_data_out3[11] .power_up = "low";

dffeas \ram_data_out0[11] (
	.clk(clk),
	.d(q_b_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_11),
	.prn(vcc));
defparam \ram_data_out0[11] .is_wysiwyg = "true";
defparam \ram_data_out0[11] .power_up = "low";

dffeas \ram_data_out1[11] (
	.clk(clk),
	.d(q_b_112),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_11),
	.prn(vcc));
defparam \ram_data_out1[11] .is_wysiwyg = "true";
defparam \ram_data_out1[11] .power_up = "low";

dffeas \ram_data_out2[10] (
	.clk(clk),
	.d(q_b_103),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_10),
	.prn(vcc));
defparam \ram_data_out2[10] .is_wysiwyg = "true";
defparam \ram_data_out2[10] .power_up = "low";

dffeas \ram_data_out3[10] (
	.clk(clk),
	.d(q_b_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_10),
	.prn(vcc));
defparam \ram_data_out3[10] .is_wysiwyg = "true";
defparam \ram_data_out3[10] .power_up = "low";

dffeas \ram_data_out0[10] (
	.clk(clk),
	.d(q_b_101),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_10),
	.prn(vcc));
defparam \ram_data_out0[10] .is_wysiwyg = "true";
defparam \ram_data_out0[10] .power_up = "low";

dffeas \ram_data_out1[10] (
	.clk(clk),
	.d(q_b_102),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_10),
	.prn(vcc));
defparam \ram_data_out1[10] .is_wysiwyg = "true";
defparam \ram_data_out1[10] .power_up = "low";

dffeas \ram_data_out0[19] (
	.clk(clk),
	.d(q_b_191),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_19),
	.prn(vcc));
defparam \ram_data_out0[19] .is_wysiwyg = "true";
defparam \ram_data_out0[19] .power_up = "low";

dffeas \ram_data_out1[19] (
	.clk(clk),
	.d(q_b_192),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_19),
	.prn(vcc));
defparam \ram_data_out1[19] .is_wysiwyg = "true";
defparam \ram_data_out1[19] .power_up = "low";

dffeas \ram_data_out2[19] (
	.clk(clk),
	.d(q_b_193),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_19),
	.prn(vcc));
defparam \ram_data_out2[19] .is_wysiwyg = "true";
defparam \ram_data_out2[19] .power_up = "low";

dffeas \ram_data_out3[19] (
	.clk(clk),
	.d(q_b_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_19),
	.prn(vcc));
defparam \ram_data_out3[19] .is_wysiwyg = "true";
defparam \ram_data_out3[19] .power_up = "low";

dffeas \ram_data_out0[5] (
	.clk(clk),
	.d(q_b_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_5),
	.prn(vcc));
defparam \ram_data_out0[5] .is_wysiwyg = "true";
defparam \ram_data_out0[5] .power_up = "low";

dffeas \ram_data_out1[5] (
	.clk(clk),
	.d(q_b_52),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_5),
	.prn(vcc));
defparam \ram_data_out1[5] .is_wysiwyg = "true";
defparam \ram_data_out1[5] .power_up = "low";

dffeas \ram_data_out2[5] (
	.clk(clk),
	.d(q_b_53),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_5),
	.prn(vcc));
defparam \ram_data_out2[5] .is_wysiwyg = "true";
defparam \ram_data_out2[5] .power_up = "low";

dffeas \ram_data_out3[5] (
	.clk(clk),
	.d(q_b_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_5),
	.prn(vcc));
defparam \ram_data_out3[5] .is_wysiwyg = "true";
defparam \ram_data_out3[5] .power_up = "low";

dffeas \ram_data_out0[6] (
	.clk(clk),
	.d(q_b_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_6),
	.prn(vcc));
defparam \ram_data_out0[6] .is_wysiwyg = "true";
defparam \ram_data_out0[6] .power_up = "low";

dffeas \ram_data_out1[6] (
	.clk(clk),
	.d(q_b_62),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_6),
	.prn(vcc));
defparam \ram_data_out1[6] .is_wysiwyg = "true";
defparam \ram_data_out1[6] .power_up = "low";

dffeas \ram_data_out2[6] (
	.clk(clk),
	.d(q_b_63),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_6),
	.prn(vcc));
defparam \ram_data_out2[6] .is_wysiwyg = "true";
defparam \ram_data_out2[6] .power_up = "low";

dffeas \ram_data_out3[6] (
	.clk(clk),
	.d(q_b_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_6),
	.prn(vcc));
defparam \ram_data_out3[6] .is_wysiwyg = "true";
defparam \ram_data_out3[6] .power_up = "low";

dffeas \ram_data_out0[7] (
	.clk(clk),
	.d(q_b_71),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_7),
	.prn(vcc));
defparam \ram_data_out0[7] .is_wysiwyg = "true";
defparam \ram_data_out0[7] .power_up = "low";

dffeas \ram_data_out1[7] (
	.clk(clk),
	.d(q_b_72),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_7),
	.prn(vcc));
defparam \ram_data_out1[7] .is_wysiwyg = "true";
defparam \ram_data_out1[7] .power_up = "low";

dffeas \ram_data_out2[7] (
	.clk(clk),
	.d(q_b_73),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_7),
	.prn(vcc));
defparam \ram_data_out2[7] .is_wysiwyg = "true";
defparam \ram_data_out2[7] .power_up = "low";

dffeas \ram_data_out3[7] (
	.clk(clk),
	.d(q_b_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_7),
	.prn(vcc));
defparam \ram_data_out3[7] .is_wysiwyg = "true";
defparam \ram_data_out3[7] .power_up = "low";

dffeas \ram_data_out0[8] (
	.clk(clk),
	.d(q_b_81),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_8),
	.prn(vcc));
defparam \ram_data_out0[8] .is_wysiwyg = "true";
defparam \ram_data_out0[8] .power_up = "low";

dffeas \ram_data_out1[8] (
	.clk(clk),
	.d(q_b_82),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_8),
	.prn(vcc));
defparam \ram_data_out1[8] .is_wysiwyg = "true";
defparam \ram_data_out1[8] .power_up = "low";

dffeas \ram_data_out2[8] (
	.clk(clk),
	.d(q_b_83),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_8),
	.prn(vcc));
defparam \ram_data_out2[8] .is_wysiwyg = "true";
defparam \ram_data_out2[8] .power_up = "low";

dffeas \ram_data_out3[8] (
	.clk(clk),
	.d(q_b_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_8),
	.prn(vcc));
defparam \ram_data_out3[8] .is_wysiwyg = "true";
defparam \ram_data_out3[8] .power_up = "low";

dffeas \ram_data_out0[4] (
	.clk(clk),
	.d(q_b_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_4),
	.prn(vcc));
defparam \ram_data_out0[4] .is_wysiwyg = "true";
defparam \ram_data_out0[4] .power_up = "low";

dffeas \ram_data_out1[4] (
	.clk(clk),
	.d(q_b_42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_4),
	.prn(vcc));
defparam \ram_data_out1[4] .is_wysiwyg = "true";
defparam \ram_data_out1[4] .power_up = "low";

dffeas \ram_data_out2[4] (
	.clk(clk),
	.d(q_b_43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_4),
	.prn(vcc));
defparam \ram_data_out2[4] .is_wysiwyg = "true";
defparam \ram_data_out2[4] .power_up = "low";

dffeas \ram_data_out3[4] (
	.clk(clk),
	.d(q_b_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_4),
	.prn(vcc));
defparam \ram_data_out3[4] .is_wysiwyg = "true";
defparam \ram_data_out3[4] .power_up = "low";

dffeas \ram_data_out2[3] (
	.clk(clk),
	.d(q_b_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_3),
	.prn(vcc));
defparam \ram_data_out2[3] .is_wysiwyg = "true";
defparam \ram_data_out2[3] .power_up = "low";

dffeas \ram_data_out3[3] (
	.clk(clk),
	.d(q_b_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_3),
	.prn(vcc));
defparam \ram_data_out3[3] .is_wysiwyg = "true";
defparam \ram_data_out3[3] .power_up = "low";

dffeas \ram_data_out0[3] (
	.clk(clk),
	.d(q_b_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_3),
	.prn(vcc));
defparam \ram_data_out0[3] .is_wysiwyg = "true";
defparam \ram_data_out0[3] .power_up = "low";

dffeas \ram_data_out1[3] (
	.clk(clk),
	.d(q_b_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_3),
	.prn(vcc));
defparam \ram_data_out1[3] .is_wysiwyg = "true";
defparam \ram_data_out1[3] .power_up = "low";

dffeas \ram_data_out2[2] (
	.clk(clk),
	.d(q_b_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_2),
	.prn(vcc));
defparam \ram_data_out2[2] .is_wysiwyg = "true";
defparam \ram_data_out2[2] .power_up = "low";

dffeas \ram_data_out3[2] (
	.clk(clk),
	.d(q_b_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_2),
	.prn(vcc));
defparam \ram_data_out3[2] .is_wysiwyg = "true";
defparam \ram_data_out3[2] .power_up = "low";

dffeas \ram_data_out0[2] (
	.clk(clk),
	.d(q_b_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_2),
	.prn(vcc));
defparam \ram_data_out0[2] .is_wysiwyg = "true";
defparam \ram_data_out0[2] .power_up = "low";

dffeas \ram_data_out1[2] (
	.clk(clk),
	.d(q_b_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_2),
	.prn(vcc));
defparam \ram_data_out1[2] .is_wysiwyg = "true";
defparam \ram_data_out1[2] .power_up = "low";

dffeas \ram_data_out2[1] (
	.clk(clk),
	.d(q_b_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_1),
	.prn(vcc));
defparam \ram_data_out2[1] .is_wysiwyg = "true";
defparam \ram_data_out2[1] .power_up = "low";

dffeas \ram_data_out3[1] (
	.clk(clk),
	.d(q_b_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_1),
	.prn(vcc));
defparam \ram_data_out3[1] .is_wysiwyg = "true";
defparam \ram_data_out3[1] .power_up = "low";

dffeas \ram_data_out0[1] (
	.clk(clk),
	.d(q_b_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_1),
	.prn(vcc));
defparam \ram_data_out0[1] .is_wysiwyg = "true";
defparam \ram_data_out0[1] .power_up = "low";

dffeas \ram_data_out1[1] (
	.clk(clk),
	.d(q_b_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_1),
	.prn(vcc));
defparam \ram_data_out1[1] .is_wysiwyg = "true";
defparam \ram_data_out1[1] .power_up = "low";

dffeas \ram_data_out2[0] (
	.clk(clk),
	.d(q_b_03),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_0),
	.prn(vcc));
defparam \ram_data_out2[0] .is_wysiwyg = "true";
defparam \ram_data_out2[0] .power_up = "low";

dffeas \ram_data_out3[0] (
	.clk(clk),
	.d(q_b_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_0),
	.prn(vcc));
defparam \ram_data_out3[0] .is_wysiwyg = "true";
defparam \ram_data_out3[0] .power_up = "low";

dffeas \ram_data_out0[0] (
	.clk(clk),
	.d(q_b_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_0),
	.prn(vcc));
defparam \ram_data_out0[0] .is_wysiwyg = "true";
defparam \ram_data_out0[0] .power_up = "low";

dffeas \ram_data_out1[0] (
	.clk(clk),
	.d(q_b_02),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_0),
	.prn(vcc));
defparam \ram_data_out1[0] .is_wysiwyg = "true";
defparam \ram_data_out1[0] .power_up = "low";

dffeas \ram_data_out0[9] (
	.clk(clk),
	.d(q_b_91),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out0_9),
	.prn(vcc));
defparam \ram_data_out0[9] .is_wysiwyg = "true";
defparam \ram_data_out0[9] .power_up = "low";

dffeas \ram_data_out1[9] (
	.clk(clk),
	.d(q_b_92),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out1_9),
	.prn(vcc));
defparam \ram_data_out1[9] .is_wysiwyg = "true";
defparam \ram_data_out1[9] .power_up = "low";

dffeas \ram_data_out2[9] (
	.clk(clk),
	.d(q_b_93),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out2_9),
	.prn(vcc));
defparam \ram_data_out2[9] .is_wysiwyg = "true";
defparam \ram_data_out2[9] .power_up = "low";

dffeas \ram_data_out3[9] (
	.clk(clk),
	.d(q_b_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(ram_data_out3_9),
	.prn(vcc));
defparam \ram_data_out3[9] .is_wysiwyg = "true";
defparam \ram_data_out3[9] .power_up = "low";

cycloneive_lcell_comb \a_ram_data_in_bus~0 (
	.dataa(ram_in_reg_2_3),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~0_combout ),
	.cout());
defparam \a_ram_data_in_bus~0 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~0 (
	.dataa(ram_in_reg_0_11),
	.datab(wr_address_i_int_0),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~0_combout ),
	.cout());
defparam \wraddress_a_bus~0 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~1 (
	.dataa(ram_in_reg_1_3),
	.datab(wr_address_i_int_1),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~1_combout ),
	.cout());
defparam \wraddress_a_bus~1 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~2 (
	.dataa(ram_in_reg_2_11),
	.datab(wr_address_i_int_2),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~2_combout ),
	.cout());
defparam \wraddress_a_bus~2 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~3 (
	.dataa(ram_in_reg_3_3),
	.datab(wr_address_i_int_3),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~3_combout ),
	.cout());
defparam \wraddress_a_bus~3 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~4 (
	.dataa(ram_in_reg_4_11),
	.datab(wr_address_i_int_4),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~4_combout ),
	.cout());
defparam \wraddress_a_bus~4 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~5 (
	.dataa(ram_in_reg_5_3),
	.datab(wr_address_i_int_5),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~5_combout ),
	.cout());
defparam \wraddress_a_bus~5 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~6 (
	.dataa(ram_block3a0),
	.datab(wr_address_i_int_6),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~6_combout ),
	.cout());
defparam \wraddress_a_bus~6 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~7 (
	.dataa(ram_block3a1),
	.datab(wr_address_i_int_7),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~7_combout ),
	.cout());
defparam \wraddress_a_bus~7 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~0 (
	.dataa(ram_in_reg_0_12),
	.datab(ram_in_reg_0_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~0_combout ),
	.cout());
defparam \rdaddress_a_bus~0 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~1 (
	.dataa(ram_in_reg_1_32),
	.datab(ram_in_reg_1_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~1_combout ),
	.cout());
defparam \rdaddress_a_bus~1 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~2 (
	.dataa(ram_in_reg_2_12),
	.datab(ram_in_reg_2_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~2_combout ),
	.cout());
defparam \rdaddress_a_bus~2 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~3 (
	.dataa(ram_in_reg_3_32),
	.datab(ram_in_reg_3_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~3_combout ),
	.cout());
defparam \rdaddress_a_bus~3 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~4 (
	.dataa(ram_in_reg_4_12),
	.datab(ram_in_reg_4_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~4_combout ),
	.cout());
defparam \rdaddress_a_bus~4 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~5 (
	.dataa(ram_in_reg_5_32),
	.datab(ram_in_reg_5_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~5_combout ),
	.cout());
defparam \rdaddress_a_bus~5 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~6 (
	.dataa(ram_in_reg_6_01),
	.datab(ram_in_reg_6_11),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~6_combout ),
	.cout());
defparam \rdaddress_a_bus~6 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~7 (
	.dataa(ram_in_reg_7_01),
	.datab(ram_in_reg_7_31),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~7_combout ),
	.cout());
defparam \rdaddress_a_bus~7 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~1 (
	.dataa(ram_in_reg_2_0),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~1_combout ),
	.cout());
defparam \a_ram_data_in_bus~1 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~8 (
	.dataa(ram_in_reg_0_02),
	.datab(wr_address_i_int_0),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~8_combout ),
	.cout());
defparam \wraddress_a_bus~8 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~9 (
	.dataa(ram_in_reg_1_0),
	.datab(wr_address_i_int_1),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~9_combout ),
	.cout());
defparam \wraddress_a_bus~9 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~10 (
	.dataa(ram_in_reg_2_02),
	.datab(wr_address_i_int_2),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~10_combout ),
	.cout());
defparam \wraddress_a_bus~10 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~11 (
	.dataa(ram_in_reg_3_0),
	.datab(wr_address_i_int_3),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~11_combout ),
	.cout());
defparam \wraddress_a_bus~11 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~12 (
	.dataa(ram_in_reg_4_02),
	.datab(wr_address_i_int_4),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~12_combout ),
	.cout());
defparam \wraddress_a_bus~12 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~13 (
	.dataa(ram_in_reg_5_0),
	.datab(wr_address_i_int_5),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~13_combout ),
	.cout());
defparam \wraddress_a_bus~13 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~8 (
	.dataa(ram_in_reg_0_03),
	.datab(ram_in_reg_0_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~8_combout ),
	.cout());
defparam \rdaddress_a_bus~8 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~9 (
	.dataa(ram_in_reg_1_03),
	.datab(ram_in_reg_1_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~9_combout ),
	.cout());
defparam \rdaddress_a_bus~9 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~10 (
	.dataa(ram_in_reg_2_03),
	.datab(ram_in_reg_2_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~10_combout ),
	.cout());
defparam \rdaddress_a_bus~10 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~11 (
	.dataa(ram_in_reg_3_03),
	.datab(ram_in_reg_3_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~11_combout ),
	.cout());
defparam \rdaddress_a_bus~11 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~12 (
	.dataa(ram_in_reg_4_03),
	.datab(ram_in_reg_4_01),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~12_combout ),
	.cout());
defparam \rdaddress_a_bus~12 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~13 (
	.dataa(ram_in_reg_5_03),
	.datab(ram_in_reg_5_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~13_combout ),
	.cout());
defparam \rdaddress_a_bus~13 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~14 (
	.dataa(ram_in_reg_6_01),
	.datab(data_rdy_vec_0),
	.datac(lpp_c_i),
	.datad(ram_in_reg_6_11),
	.cin(gnd),
	.combout(\rdaddress_a_bus~14_combout ),
	.cout());
defparam \rdaddress_a_bus~14 .lut_mask = 16'hBEFF;
defparam \rdaddress_a_bus~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~15 (
	.dataa(ram_in_reg_7_01),
	.datab(data_rdy_vec_0),
	.datac(lpp_c_i),
	.datad(ram_in_reg_7_21),
	.cin(gnd),
	.combout(\rdaddress_a_bus~15_combout ),
	.cout());
defparam \rdaddress_a_bus~15 .lut_mask = 16'hBEFF;
defparam \rdaddress_a_bus~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~2 (
	.dataa(ram_in_reg_2_1),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~2_combout ),
	.cout());
defparam \a_ram_data_in_bus~2 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~14 (
	.dataa(ram_in_reg_1_1),
	.datab(wr_address_i_int_1),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~14_combout ),
	.cout());
defparam \wraddress_a_bus~14 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~15 (
	.dataa(ram_in_reg_3_1),
	.datab(wr_address_i_int_3),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~15_combout ),
	.cout());
defparam \wraddress_a_bus~15 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~16 (
	.dataa(ram_in_reg_5_1),
	.datab(wr_address_i_int_5),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~16_combout ),
	.cout());
defparam \wraddress_a_bus~16 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~16 (
	.dataa(ram_in_reg_1_12),
	.datab(ram_in_reg_1_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~16_combout ),
	.cout());
defparam \rdaddress_a_bus~16 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~17 (
	.dataa(ram_in_reg_3_12),
	.datab(ram_in_reg_3_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~17_combout ),
	.cout());
defparam \rdaddress_a_bus~17 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~18 (
	.dataa(ram_in_reg_5_12),
	.datab(ram_in_reg_5_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~18_combout ),
	.cout());
defparam \rdaddress_a_bus~18 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~19 (
	.dataa(ram_in_reg_7_01),
	.datab(data_rdy_vec_0),
	.datac(lpp_c_i),
	.datad(ram_in_reg_7_31),
	.cin(gnd),
	.combout(\rdaddress_a_bus~19_combout ),
	.cout());
defparam \rdaddress_a_bus~19 .lut_mask = 16'hBEFF;
defparam \rdaddress_a_bus~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~3 (
	.dataa(ram_in_reg_2_2),
	.datab(data_in_r_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~3_combout ),
	.cout());
defparam \a_ram_data_in_bus~3 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~17 (
	.dataa(ram_in_reg_1_2),
	.datab(wr_address_i_int_1),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~17_combout ),
	.cout());
defparam \wraddress_a_bus~17 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~18 (
	.dataa(ram_in_reg_3_2),
	.datab(wr_address_i_int_3),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~18_combout ),
	.cout());
defparam \wraddress_a_bus~18 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wraddress_a_bus~19 (
	.dataa(ram_in_reg_5_2),
	.datab(wr_address_i_int_5),
	.datac(wc_vec_3),
	.datad(data_rdy_vec_2),
	.cin(gnd),
	.combout(\wraddress_a_bus~19_combout ),
	.cout());
defparam \wraddress_a_bus~19 .lut_mask = 16'hEFFE;
defparam \wraddress_a_bus~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~20 (
	.dataa(ram_in_reg_1_22),
	.datab(ram_in_reg_1_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~20_combout ),
	.cout());
defparam \rdaddress_a_bus~20 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~21 (
	.dataa(ram_in_reg_3_22),
	.datab(ram_in_reg_3_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~21_combout ),
	.cout());
defparam \rdaddress_a_bus~21 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~22 (
	.dataa(ram_in_reg_5_22),
	.datab(ram_in_reg_5_02),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~22_combout ),
	.cout());
defparam \rdaddress_a_bus~22 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdaddress_a_bus~23 (
	.dataa(ram_in_reg_7_01),
	.datab(ram_in_reg_7_21),
	.datac(lpp_c_i),
	.datad(data_rdy_vec_0),
	.cin(gnd),
	.combout(\rdaddress_a_bus~23_combout ),
	.cout());
defparam \rdaddress_a_bus~23 .lut_mask = 16'hEFFE;
defparam \rdaddress_a_bus~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~4 (
	.dataa(ram_in_reg_2_7),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~4_combout ),
	.cout());
defparam \a_ram_data_in_bus~4 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~5 (
	.dataa(ram_in_reg_2_4),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~5_combout ),
	.cout());
defparam \a_ram_data_in_bus~5 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~6 (
	.dataa(ram_in_reg_2_5),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~6_combout ),
	.cout());
defparam \a_ram_data_in_bus~6 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~7 (
	.dataa(ram_in_reg_2_6),
	.datab(data_in_i_2),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~7_combout ),
	.cout());
defparam \a_ram_data_in_bus~7 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~8 (
	.dataa(ram_in_reg_1_31),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~8_combout ),
	.cout());
defparam \a_ram_data_in_bus~8 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~9 (
	.dataa(ram_in_reg_1_01),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~9_combout ),
	.cout());
defparam \a_ram_data_in_bus~9 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~10 (
	.dataa(ram_in_reg_1_11),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~10_combout ),
	.cout());
defparam \a_ram_data_in_bus~10 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~11 (
	.dataa(ram_in_reg_1_21),
	.datab(data_in_r_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~11_combout ),
	.cout());
defparam \a_ram_data_in_bus~11 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~12 (
	.dataa(ram_in_reg_1_7),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~12_combout ),
	.cout());
defparam \a_ram_data_in_bus~12 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~13 (
	.dataa(ram_in_reg_1_4),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~13_combout ),
	.cout());
defparam \a_ram_data_in_bus~13 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~14 (
	.dataa(ram_in_reg_1_5),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~14_combout ),
	.cout());
defparam \a_ram_data_in_bus~14 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~15 (
	.dataa(ram_in_reg_1_6),
	.datab(data_in_i_1),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~15_combout ),
	.cout());
defparam \a_ram_data_in_bus~15 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~16 (
	.dataa(ram_in_reg_0_3),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~16_combout ),
	.cout());
defparam \a_ram_data_in_bus~16 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~17 (
	.dataa(ram_in_reg_0_0),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~17_combout ),
	.cout());
defparam \a_ram_data_in_bus~17 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~18 (
	.dataa(ram_in_reg_0_1),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~18_combout ),
	.cout());
defparam \a_ram_data_in_bus~18 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~19 (
	.dataa(ram_in_reg_0_2),
	.datab(data_in_r_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~19_combout ),
	.cout());
defparam \a_ram_data_in_bus~19 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~20 (
	.dataa(ram_in_reg_0_7),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~20_combout ),
	.cout());
defparam \a_ram_data_in_bus~20 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~21 (
	.dataa(ram_in_reg_0_4),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~21_combout ),
	.cout());
defparam \a_ram_data_in_bus~21 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~22 (
	.dataa(ram_in_reg_0_5),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~22_combout ),
	.cout());
defparam \a_ram_data_in_bus~22 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~23 (
	.dataa(ram_in_reg_0_6),
	.datab(data_in_i_0),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~23_combout ),
	.cout());
defparam \a_ram_data_in_bus~23 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~24 (
	.dataa(ram_in_reg_9_3),
	.datab(data_in_r_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~24_combout ),
	.cout());
defparam \a_ram_data_in_bus~24 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~25 (
	.dataa(ram_in_reg_9_0),
	.datab(data_in_r_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~25_combout ),
	.cout());
defparam \a_ram_data_in_bus~25 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~26 (
	.dataa(ram_in_reg_9_1),
	.datab(data_in_r_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~26_combout ),
	.cout());
defparam \a_ram_data_in_bus~26 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~27 (
	.dataa(ram_in_reg_9_2),
	.datab(data_in_r_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~27_combout ),
	.cout());
defparam \a_ram_data_in_bus~27 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~28 (
	.dataa(ram_in_reg_9_7),
	.datab(data_in_i_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~28_combout ),
	.cout());
defparam \a_ram_data_in_bus~28 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~29 (
	.dataa(ram_in_reg_9_4),
	.datab(data_in_i_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~29_combout ),
	.cout());
defparam \a_ram_data_in_bus~29 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~30 (
	.dataa(ram_in_reg_9_5),
	.datab(data_in_i_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~30_combout ),
	.cout());
defparam \a_ram_data_in_bus~30 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~31 (
	.dataa(ram_in_reg_9_6),
	.datab(data_in_i_9),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~31_combout ),
	.cout());
defparam \a_ram_data_in_bus~31 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~32 (
	.dataa(ram_in_reg_8_3),
	.datab(data_in_r_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~32_combout ),
	.cout());
defparam \a_ram_data_in_bus~32 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~33 (
	.dataa(ram_in_reg_8_0),
	.datab(data_in_r_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~33_combout ),
	.cout());
defparam \a_ram_data_in_bus~33 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~34 (
	.dataa(ram_in_reg_8_1),
	.datab(data_in_r_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~34_combout ),
	.cout());
defparam \a_ram_data_in_bus~34 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~35 (
	.dataa(ram_in_reg_8_2),
	.datab(data_in_r_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~35_combout ),
	.cout());
defparam \a_ram_data_in_bus~35 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~36 (
	.dataa(ram_in_reg_8_7),
	.datab(data_in_i_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~36_combout ),
	.cout());
defparam \a_ram_data_in_bus~36 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~37 (
	.dataa(ram_in_reg_8_4),
	.datab(data_in_i_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~37_combout ),
	.cout());
defparam \a_ram_data_in_bus~37 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~38 (
	.dataa(ram_in_reg_8_5),
	.datab(data_in_i_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~38_combout ),
	.cout());
defparam \a_ram_data_in_bus~38 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~39 (
	.dataa(ram_in_reg_8_6),
	.datab(data_in_i_8),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~39_combout ),
	.cout());
defparam \a_ram_data_in_bus~39 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~40 (
	.dataa(ram_in_reg_7_3),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~40_combout ),
	.cout());
defparam \a_ram_data_in_bus~40 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~41 (
	.dataa(ram_in_reg_7_0),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~41_combout ),
	.cout());
defparam \a_ram_data_in_bus~41 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~42 (
	.dataa(ram_in_reg_7_1),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~42_combout ),
	.cout());
defparam \a_ram_data_in_bus~42 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~43 (
	.dataa(ram_in_reg_7_2),
	.datab(data_in_r_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~43_combout ),
	.cout());
defparam \a_ram_data_in_bus~43 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~44 (
	.dataa(ram_in_reg_7_7),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~44_combout ),
	.cout());
defparam \a_ram_data_in_bus~44 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~45 (
	.dataa(ram_in_reg_7_4),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~45_combout ),
	.cout());
defparam \a_ram_data_in_bus~45 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~46 (
	.dataa(ram_in_reg_7_5),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~46_combout ),
	.cout());
defparam \a_ram_data_in_bus~46 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~47 (
	.dataa(ram_in_reg_7_6),
	.datab(data_in_i_7),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~47_combout ),
	.cout());
defparam \a_ram_data_in_bus~47 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~48 (
	.dataa(ram_in_reg_6_3),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~48_combout ),
	.cout());
defparam \a_ram_data_in_bus~48 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~49 (
	.dataa(ram_in_reg_6_0),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~49_combout ),
	.cout());
defparam \a_ram_data_in_bus~49 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~50 (
	.dataa(ram_in_reg_6_1),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~50_combout ),
	.cout());
defparam \a_ram_data_in_bus~50 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~51 (
	.dataa(ram_in_reg_6_2),
	.datab(data_in_r_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~51_combout ),
	.cout());
defparam \a_ram_data_in_bus~51 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~52 (
	.dataa(ram_in_reg_6_7),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~52_combout ),
	.cout());
defparam \a_ram_data_in_bus~52 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~53 (
	.dataa(ram_in_reg_6_4),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~53_combout ),
	.cout());
defparam \a_ram_data_in_bus~53 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~54 (
	.dataa(ram_in_reg_6_5),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~54_combout ),
	.cout());
defparam \a_ram_data_in_bus~54 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~55 (
	.dataa(ram_in_reg_6_6),
	.datab(data_in_i_6),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~55_combout ),
	.cout());
defparam \a_ram_data_in_bus~55 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~56 (
	.dataa(ram_in_reg_5_31),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~56_combout ),
	.cout());
defparam \a_ram_data_in_bus~56 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~57 (
	.dataa(ram_in_reg_5_01),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~57_combout ),
	.cout());
defparam \a_ram_data_in_bus~57 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~58 (
	.dataa(ram_in_reg_5_11),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~58_combout ),
	.cout());
defparam \a_ram_data_in_bus~58 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~59 (
	.dataa(ram_in_reg_5_21),
	.datab(data_in_r_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~59_combout ),
	.cout());
defparam \a_ram_data_in_bus~59 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~60 (
	.dataa(ram_in_reg_5_7),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~60_combout ),
	.cout());
defparam \a_ram_data_in_bus~60 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~61 (
	.dataa(ram_in_reg_5_4),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~61_combout ),
	.cout());
defparam \a_ram_data_in_bus~61 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~62 (
	.dataa(ram_in_reg_5_5),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~62_combout ),
	.cout());
defparam \a_ram_data_in_bus~62 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~63 (
	.dataa(ram_in_reg_5_6),
	.datab(data_in_i_5),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~63_combout ),
	.cout());
defparam \a_ram_data_in_bus~63 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~64 (
	.dataa(ram_in_reg_4_3),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~64_combout ),
	.cout());
defparam \a_ram_data_in_bus~64 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~65 (
	.dataa(ram_in_reg_4_0),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~65_combout ),
	.cout());
defparam \a_ram_data_in_bus~65 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~66 (
	.dataa(ram_in_reg_4_1),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~66_combout ),
	.cout());
defparam \a_ram_data_in_bus~66 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~67 (
	.dataa(ram_in_reg_4_2),
	.datab(data_in_r_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~67_combout ),
	.cout());
defparam \a_ram_data_in_bus~67 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~68 (
	.dataa(ram_in_reg_4_7),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~68_combout ),
	.cout());
defparam \a_ram_data_in_bus~68 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~69 (
	.dataa(ram_in_reg_4_4),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~69_combout ),
	.cout());
defparam \a_ram_data_in_bus~69 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~70 (
	.dataa(ram_in_reg_4_5),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~70_combout ),
	.cout());
defparam \a_ram_data_in_bus~70 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~71 (
	.dataa(ram_in_reg_4_6),
	.datab(data_in_i_4),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~71_combout ),
	.cout());
defparam \a_ram_data_in_bus~71 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~72 (
	.dataa(ram_in_reg_3_31),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~72_combout ),
	.cout());
defparam \a_ram_data_in_bus~72 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~73 (
	.dataa(ram_in_reg_3_01),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~73_combout ),
	.cout());
defparam \a_ram_data_in_bus~73 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~74 (
	.dataa(ram_in_reg_3_11),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~74_combout ),
	.cout());
defparam \a_ram_data_in_bus~74 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~75 (
	.dataa(ram_in_reg_3_21),
	.datab(data_in_r_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~75_combout ),
	.cout());
defparam \a_ram_data_in_bus~75 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~76 (
	.dataa(ram_in_reg_3_7),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~76_combout ),
	.cout());
defparam \a_ram_data_in_bus~76 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~77 (
	.dataa(ram_in_reg_3_4),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~77_combout ),
	.cout());
defparam \a_ram_data_in_bus~77 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~78 (
	.dataa(ram_in_reg_3_5),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~78_combout ),
	.cout());
defparam \a_ram_data_in_bus~78 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \a_ram_data_in_bus~79 (
	.dataa(ram_in_reg_3_6),
	.datab(data_in_i_3),
	.datac(gnd),
	.datad(sel_ram_in),
	.cin(gnd),
	.combout(\a_ram_data_in_bus~79_combout ),
	.cout());
defparam \a_ram_data_in_bus~79 .lut_mask = 16'hAACC;
defparam \a_ram_data_in_bus~79 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_wrengen (
	lpp_c_i1,
	global_clock_enable,
	stall_reg,
	source_stall_int_d,
	global_clock_enable1,
	wait_count_0,
	wc_i_d1,
	p_cd_en_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	lpp_c_i1;
input 	global_clock_enable;
input 	stall_reg;
input 	source_stall_int_d;
input 	global_clock_enable1;
output 	wait_count_0;
output 	wc_i_d1;
input 	p_cd_en_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wc_state.IDLE~0_combout ;
wire \wc_state.IDLE~q ;
wire \wait_count~3_combout ;
wire \wait_count[0]~q ;
wire \wait_count~4_combout ;
wire \wait_count[1]~q ;
wire \wait_count~1_combout ;
wire \wait_count[2]~q ;
wire \Add0~0_combout ;
wire \wait_count~2_combout ;
wire \wait_count[3]~q ;
wire \Selector2~0_combout ;
wire \Selector1~0_combout ;
wire \wc_state.WAIT_LAT~q ;
wire \Selector2~1_combout ;
wire \wc_state.ENABLE~q ;
wire \wc_i~q ;
wire \lpp_c_i~0_combout ;
wire \wc_i_d~0_combout ;


dffeas lpp_c_i(
	.clk(clk),
	.d(\lpp_c_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(lpp_c_i1),
	.prn(vcc));
defparam lpp_c_i.is_wysiwyg = "true";
defparam lpp_c_i.power_up = "low";

cycloneive_lcell_comb \wait_count[0]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(global_clock_enable),
	.datad(source_stall_int_d),
	.cin(gnd),
	.combout(wait_count_0),
	.cout());
defparam \wait_count[0]~0 .lut_mask = 16'hACFF;
defparam \wait_count[0]~0 .sum_lutc_input = "datac";

dffeas wc_i_d(
	.clk(clk),
	.d(\wc_i_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(wc_i_d1),
	.prn(vcc));
defparam wc_i_d.is_wysiwyg = "true";
defparam wc_i_d.power_up = "low";

cycloneive_lcell_comb \wc_state.IDLE~0 (
	.dataa(gnd),
	.datab(p_cd_en_2),
	.datac(\wc_state.WAIT_LAT~q ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\wc_state.IDLE~0_combout ),
	.cout());
defparam \wc_state.IDLE~0 .lut_mask = 16'hFFFC;
defparam \wc_state.IDLE~0 .sum_lutc_input = "datac";

dffeas \wc_state.IDLE (
	.clk(clk),
	.d(\wc_state.IDLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(\wc_state.IDLE~q ),
	.prn(vcc));
defparam \wc_state.IDLE .is_wysiwyg = "true";
defparam \wc_state.IDLE .power_up = "low";

cycloneive_lcell_comb \wait_count~3 (
	.dataa(\wait_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wc_state.WAIT_LAT~q ),
	.cin(gnd),
	.combout(\wait_count~3_combout ),
	.cout());
defparam \wait_count~3 .lut_mask = 16'hFF55;
defparam \wait_count~3 .sum_lutc_input = "datac";

dffeas \wait_count[0] (
	.clk(clk),
	.d(\wait_count~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(\wait_count[0]~q ),
	.prn(vcc));
defparam \wait_count[0] .is_wysiwyg = "true";
defparam \wait_count[0] .power_up = "low";

cycloneive_lcell_comb \wait_count~4 (
	.dataa(\wc_state.WAIT_LAT~q ),
	.datab(gnd),
	.datac(\wait_count[0]~q ),
	.datad(\wait_count[1]~q ),
	.cin(gnd),
	.combout(\wait_count~4_combout ),
	.cout());
defparam \wait_count~4 .lut_mask = 16'hAFFA;
defparam \wait_count~4 .sum_lutc_input = "datac";

dffeas \wait_count[1] (
	.clk(clk),
	.d(\wait_count~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(\wait_count[1]~q ),
	.prn(vcc));
defparam \wait_count[1] .is_wysiwyg = "true";
defparam \wait_count[1] .power_up = "low";

cycloneive_lcell_comb \wait_count~1 (
	.dataa(\wc_state.WAIT_LAT~q ),
	.datab(\wait_count[2]~q ),
	.datac(\wait_count[0]~q ),
	.datad(\wait_count[1]~q ),
	.cin(gnd),
	.combout(\wait_count~1_combout ),
	.cout());
defparam \wait_count~1 .lut_mask = 16'hEBBE;
defparam \wait_count~1 .sum_lutc_input = "datac";

dffeas \wait_count[2] (
	.clk(clk),
	.d(\wait_count~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(\wait_count[2]~q ),
	.prn(vcc));
defparam \wait_count[2] .is_wysiwyg = "true";
defparam \wait_count[2] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\wait_count[3]~q ),
	.datab(\wait_count[0]~q ),
	.datac(\wait_count[1]~q ),
	.datad(\wait_count[2]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h6996;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_count~2 (
	.dataa(\wc_state.WAIT_LAT~q ),
	.datab(\Add0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wait_count~2_combout ),
	.cout());
defparam \wait_count~2 .lut_mask = 16'hEEEE;
defparam \wait_count~2 .sum_lutc_input = "datac";

dffeas \wait_count[3] (
	.clk(clk),
	.d(\wait_count~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wait_count_0),
	.q(\wait_count[3]~q ),
	.prn(vcc));
defparam \wait_count[3] .is_wysiwyg = "true";
defparam \wait_count[3] .power_up = "low";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\wait_count[2]~q ),
	.datab(\wait_count[3]~q ),
	.datac(\wait_count[0]~q ),
	.datad(\wait_count[1]~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEFFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(p_cd_en_2),
	.datab(\wc_state.WAIT_LAT~q ),
	.datac(\wc_state.IDLE~q ),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hEFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \wc_state.WAIT_LAT (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(\wc_state.WAIT_LAT~q ),
	.prn(vcc));
defparam \wc_state.WAIT_LAT .is_wysiwyg = "true";
defparam \wc_state.WAIT_LAT .power_up = "low";

cycloneive_lcell_comb \Selector2~1 (
	.dataa(\wc_state.ENABLE~q ),
	.datab(\wc_state.WAIT_LAT~q ),
	.datac(\Selector2~0_combout ),
	.datad(p_cd_en_2),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFFFE;
defparam \Selector2~1 .sum_lutc_input = "datac";

dffeas \wc_state.ENABLE (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(\wc_state.ENABLE~q ),
	.prn(vcc));
defparam \wc_state.ENABLE .is_wysiwyg = "true";
defparam \wc_state.ENABLE .power_up = "low";

dffeas wc_i(
	.clk(clk),
	.d(\wc_state.ENABLE~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable1),
	.q(\wc_i~q ),
	.prn(vcc));
defparam wc_i.is_wysiwyg = "true";
defparam wc_i.power_up = "low";

cycloneive_lcell_comb \lpp_c_i~0 (
	.dataa(lpp_c_i1),
	.datab(wc_i_d1),
	.datac(gnd),
	.datad(\wc_i~q ),
	.cin(gnd),
	.combout(\lpp_c_i~0_combout ),
	.cout());
defparam \lpp_c_i~0 .lut_mask = 16'hEEFF;
defparam \lpp_c_i~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wc_i_d~0 (
	.dataa(reset_n),
	.datab(\wc_i~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wc_i_d~0_combout ),
	.cout());
defparam \wc_i_d~0 .lut_mask = 16'hEEEE;
defparam \wc_i_d~0 .sum_lutc_input = "datac";

endmodule

module fftsign_asj_fft_wrswgen (
	ram_block3a1,
	ram_block3a0,
	ram_block3a2,
	ram_block3a3,
	global_clock_enable,
	swa_tdl_0_16,
	swa_tdl_1_16,
	p_2,
	p_0,
	p_1,
	Add1,
	Mux1,
	Mux11,
	k_count_6,
	Add0,
	Add11,
	Add12,
	Mux0,
	Mux01,
	k_count_7,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block3a1;
output 	ram_block3a0;
input 	ram_block3a2;
input 	ram_block3a3;
input 	global_clock_enable;
output 	swa_tdl_0_16;
output 	swa_tdl_1_16;
input 	p_2;
input 	p_0;
input 	p_1;
input 	Add1;
input 	Mux1;
input 	Mux11;
input 	k_count_6;
input 	Add0;
input 	Add11;
input 	Add12;
input 	Mux0;
input 	Mux01;
input 	k_count_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux0~0_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ;
wire \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ;
wire \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ;
wire \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \swd_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ;
wire \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \Add2~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \swa_tdl[15][0]~q ;
wire \swa_tdl[15][1]~q ;

wire [143:0] \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ;
wire [143:0] \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ;

assign ram_block3a1 = \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus [0];

assign ram_block3a0 = \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus [0];

cycloneive_ram_block \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux1~2_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swd_rtl_0|auto_generated|altsyncram2|ram_block3a1_PORTBDATAOUT_bus ));
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_core_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_input_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .clk0_output_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_offset_in_bits = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .data_interleave_width_in_bits = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_wrswgen:get_wr_swtiches|altshift_taps:swd_rtl_0|shift_taps_qnm:auto_generated|altsyncram_4e81:altsyncram2|ALTSYNCRAM";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .mixed_port_feed_through_mode = "old";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .operation_mode = "dual_port";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_address_width = 4;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_out_clock = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_data_width = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_address = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_first_bit_number = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_last_address = 15;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_depth = 16;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_logical_ram_width = 2;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_address_width = 4;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_out_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_data_width = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_address = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_first_bit_number = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_last_address = 15;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_depth = 16;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_logical_ram_width = 2;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .port_b_read_enable_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a1 .ram_block_type = "auto";

cycloneive_ram_block \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(global_clock_enable),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux0~3_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swd_rtl_0|auto_generated|altsyncram2|ram_block3a0_PORTBDATAOUT_bus ));
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_core_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_input_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .clk0_output_clock_enable = "ena0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_offset_in_bits = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .data_interleave_width_in_bits = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|asj_fft_wrswgen:get_wr_swtiches|altshift_taps:swd_rtl_0|shift_taps_qnm:auto_generated|altsyncram_4e81:altsyncram2|ALTSYNCRAM";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .mixed_port_feed_through_mode = "old";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .operation_mode = "dual_port";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_address_width = 4;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_out_clock = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_data_width = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_address = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_first_bit_number = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_last_address = 15;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_depth = 16;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_logical_ram_width = 2;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_address_width = 4;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clear = "none";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_out_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_data_width = 1;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_address = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_first_bit_number = 0;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_last_address = 15;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_depth = 16;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_logical_ram_width = 2;
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .port_b_read_enable_clock = "clock0";
defparam \swd_rtl_0|auto_generated|altsyncram2|ram_block3a0 .ram_block_type = "auto";

dffeas \swa_tdl[16][0] (
	.clk(clk),
	.d(\swa_tdl[15][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(swa_tdl_0_16),
	.prn(vcc));
defparam \swa_tdl[16][0] .is_wysiwyg = "true";
defparam \swa_tdl[16][0] .power_up = "low";

dffeas \swa_tdl[16][1] (
	.clk(clk),
	.d(\swa_tdl[15][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(swa_tdl_1_16),
	.prn(vcc));
defparam \swa_tdl[16][1] .is_wysiwyg = "true";
defparam \swa_tdl[16][1] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(p_1),
	.datab(gnd),
	.datac(p_2),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hAFFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(p_2),
	.datab(gnd),
	.datac(Add1),
	.datad(k_count_6),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hAFFA;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(Mux11),
	.datab(\Mux1~0_combout ),
	.datac(p_1),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hEFFE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(Add1),
	.datab(Mux1),
	.datac(\Mux0~0_combout ),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hEFFE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \swd_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ),
	.cout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ));
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita0 .sum_lutc_input = "cin";

dffeas \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb \swd_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.combout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ),
	.cout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ));
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita1 .sum_lutc_input = "cin";

dffeas \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb \swd_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.combout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ),
	.cout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ));
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita2 .sum_lutc_input = "cin";

dffeas \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb \swd_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.combout(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ),
	.cout());
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 16'h5A5A;
defparam \swd_rtl_0|auto_generated|cntr1|counter_comb_bita3 .sum_lutc_input = "cin";

dffeas \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\swd_rtl_0|auto_generated|cntr1|counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \swd_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(gnd),
	.datab(k_count_7),
	.datac(Add1),
	.datad(k_count_6),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'hC33C;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(p_2),
	.datab(Add0),
	.datac(Add11),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hEBBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(Mux01),
	.datab(\Mux0~1_combout ),
	.datac(p_1),
	.datad(p_0),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hEFFE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(Add12),
	.datab(Mux0),
	.datac(\Mux0~0_combout ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hEFFE;
defparam \Mux0~3 .sum_lutc_input = "datac";

dffeas \swa_tdl[15][0] (
	.clk(clk),
	.d(ram_block3a2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swa_tdl[15][0]~q ),
	.prn(vcc));
defparam \swa_tdl[15][0] .is_wysiwyg = "true";
defparam \swa_tdl[15][0] .power_up = "low";

dffeas \swa_tdl[15][1] (
	.clk(clk),
	.d(ram_block3a3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(global_clock_enable),
	.q(\swa_tdl[15][1]~q ),
	.prn(vcc));
defparam \swa_tdl[15][1] .is_wysiwyg = "true";
defparam \swa_tdl[15][1] .power_up = "low";

endmodule

module fftsign_auk_dspip_avalon_streaming_controller (
	master_sink_ena,
	sink_in_work,
	source_packet_error_1,
	source_packet_error_0,
	source_stall_reg1,
	sink_stall_reg1,
	send_eop_s,
	sink_ready_ctrl,
	sink_start,
	empty_dff,
	sink_stall,
	packet_error_s_1,
	packet_error_s_0,
	stall_reg1,
	Mux0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	master_sink_ena;
input 	sink_in_work;
output 	source_packet_error_1;
output 	source_packet_error_0;
output 	source_stall_reg1;
output 	sink_stall_reg1;
input 	send_eop_s;
output 	sink_ready_ctrl;
input 	sink_start;
input 	empty_dff;
input 	sink_stall;
input 	packet_error_s_1;
input 	packet_error_s_0;
output 	stall_reg1;
input 	Mux0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_stall_reg~0_combout ;
wire \sink_stall_reg~0_combout ;
wire \sink_ready_ctrl~0_combout ;
wire \stall_int~combout ;


dffeas \source_packet_error[1] (
	.clk(clk),
	.d(packet_error_s_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_1),
	.prn(vcc));
defparam \source_packet_error[1] .is_wysiwyg = "true";
defparam \source_packet_error[1] .power_up = "low";

dffeas \source_packet_error[0] (
	.clk(clk),
	.d(packet_error_s_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_0),
	.prn(vcc));
defparam \source_packet_error[0] .is_wysiwyg = "true";
defparam \source_packet_error[0] .power_up = "low";

dffeas source_stall_reg(
	.clk(clk),
	.d(\source_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_reg1),
	.prn(vcc));
defparam source_stall_reg.is_wysiwyg = "true";
defparam source_stall_reg.power_up = "low";

dffeas sink_stall_reg(
	.clk(clk),
	.d(\sink_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_stall_reg1),
	.prn(vcc));
defparam sink_stall_reg.is_wysiwyg = "true";
defparam sink_stall_reg.power_up = "low";

cycloneive_lcell_comb \sink_ready_ctrl~1 (
	.dataa(\sink_ready_ctrl~0_combout ),
	.datab(master_sink_ena),
	.datac(sink_in_work),
	.datad(send_eop_s),
	.cin(gnd),
	.combout(sink_ready_ctrl),
	.cout());
defparam \sink_ready_ctrl~1 .lut_mask = 16'hFEFF;
defparam \sink_ready_ctrl~1 .sum_lutc_input = "datac";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_int~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

cycloneive_lcell_comb \source_stall_reg~0 (
	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_stall_reg~0_combout ),
	.cout());
defparam \source_stall_reg~0 .lut_mask = 16'h5555;
defparam \source_stall_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_stall_reg~0 (
	.dataa(sink_stall),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_stall_reg~0_combout ),
	.cout());
defparam \sink_stall_reg~0 .lut_mask = 16'h5555;
defparam \sink_stall_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready_ctrl~0 (
	.dataa(source_stall_reg1),
	.datab(gnd),
	.datac(gnd),
	.datad(sink_stall_reg1),
	.cin(gnd),
	.combout(\sink_ready_ctrl~0_combout ),
	.cout());
defparam \sink_ready_ctrl~0 .lut_mask = 16'hAAFF;
defparam \sink_ready_ctrl~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb stall_int(
	.dataa(sink_start),
	.datab(empty_dff),
	.datac(Mux0),
	.datad(gnd),
	.cin(gnd),
	.combout(\stall_int~combout ),
	.cout());
defparam stall_int.lut_mask = 16'hEFEF;
defparam stall_int.sum_lutc_input = "datac";

endmodule

module fftsign_auk_dspip_avalon_streaming_sink (
	q_b_2,
	q_b_12,
	q_b_1,
	q_b_11,
	q_b_0,
	q_b_10,
	q_b_9,
	q_b_19,
	q_b_8,
	q_b_18,
	q_b_7,
	q_b_17,
	q_b_6,
	q_b_16,
	q_b_5,
	q_b_15,
	q_b_4,
	q_b_14,
	q_b_3,
	q_b_13,
	at_sink_ready_s1,
	send_eop_s1,
	sink_ready_ctrl,
	sink_start1,
	empty_dff,
	sink_stall1,
	packet_error_s_1,
	packet_error_s_0,
	send_sop_s1,
	clk,
	reset_n,
	sink_valid,
	sink_eop,
	sink_sop,
	sink_error_0,
	sink_error_1,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
output 	q_b_2;
output 	q_b_12;
output 	q_b_1;
output 	q_b_11;
output 	q_b_0;
output 	q_b_10;
output 	q_b_9;
output 	q_b_19;
output 	q_b_8;
output 	q_b_18;
output 	q_b_7;
output 	q_b_17;
output 	q_b_6;
output 	q_b_16;
output 	q_b_5;
output 	q_b_15;
output 	q_b_4;
output 	q_b_14;
output 	q_b_3;
output 	q_b_13;
output 	at_sink_ready_s1;
output 	send_eop_s1;
input 	sink_ready_ctrl;
output 	sink_start1;
output 	empty_dff;
output 	sink_stall1;
output 	packet_error_s_1;
output 	packet_error_s_0;
output 	send_sop_s1;
input 	clk;
input 	reset_n;
input 	sink_valid;
input 	sink_eop;
input 	sink_sop;
input 	sink_error_0;
input 	sink_error_1;
input 	[19:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ;
wire \fifo_wrreq~0_combout ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \at_sink_data_int[2]~q ;
wire \at_sink_data_int[12]~q ;
wire \at_sink_data_int[1]~q ;
wire \at_sink_data_int[11]~q ;
wire \at_sink_data_int[0]~q ;
wire \at_sink_data_int[10]~q ;
wire \at_sink_data_int[9]~q ;
wire \at_sink_data_int[19]~q ;
wire \at_sink_data_int[8]~q ;
wire \at_sink_data_int[18]~q ;
wire \at_sink_data_int[7]~q ;
wire \at_sink_data_int[17]~q ;
wire \at_sink_data_int[6]~q ;
wire \at_sink_data_int[16]~q ;
wire \at_sink_data_int[5]~q ;
wire \at_sink_data_int[15]~q ;
wire \at_sink_data_int[4]~q ;
wire \at_sink_data_int[14]~q ;
wire \at_sink_data_int[3]~q ;
wire \at_sink_data_int[13]~q ;
wire \data_take~combout ;
wire \at_sink_ready_s~0_combout ;
wire \out_cnt[0]~10_combout ;
wire \sink_stall_s~q ;
wire \Selector8~0_combout ;
wire \sink_out_state.normal~q ;
wire \Selector10~2_combout ;
wire \Selector10~3_combout ;
wire \sink_out_state.empty_and_ready~q ;
wire \Selector7~0_combout ;
wire \out_cnt[0]~q ;
wire \out_cnt[0]~11 ;
wire \out_cnt[1]~12_combout ;
wire \out_cnt[1]~q ;
wire \out_cnt[1]~13 ;
wire \out_cnt[2]~14_combout ;
wire \out_cnt[2]~q ;
wire \out_cnt[2]~15 ;
wire \out_cnt[3]~16_combout ;
wire \out_cnt[3]~q ;
wire \Equal2~0_combout ;
wire \out_cnt[3]~17 ;
wire \out_cnt[4]~18_combout ;
wire \out_cnt[4]~q ;
wire \out_cnt[4]~19 ;
wire \out_cnt[5]~20_combout ;
wire \out_cnt[5]~q ;
wire \out_cnt[5]~21 ;
wire \out_cnt[6]~22_combout ;
wire \out_cnt[6]~q ;
wire \out_cnt[6]~23 ;
wire \out_cnt[7]~24_combout ;
wire \out_cnt[7]~q ;
wire \Equal2~1_combout ;
wire \out_cnt[7]~25 ;
wire \out_cnt[8]~26_combout ;
wire \out_cnt[8]~q ;
wire \out_cnt[8]~27 ;
wire \out_cnt[9]~28_combout ;
wire \out_cnt[9]~q ;
wire \Equal2~2_combout ;
wire \send_sop_eop_p~0_combout ;
wire \sink_start~0_combout ;
wire \sink_comb_update_2~1_combout ;
wire \count[0]~10_combout ;
wire \Selector1~0_combout ;
wire \sink_state.stall~q ;
wire \Selector3~0_combout ;
wire \Selector2~6_combout ;
wire \Selector2~7_combout ;
wire \sink_comb_update_2~2_combout ;
wire \sink_state.st_err~q ;
wire \Selector3~2_combout ;
wire \Selector2~2_combout ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \Selector2~3_combout ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \Selector3~3_combout ;
wire \count[6]~14_combout ;
wire \Selector4~0_combout ;
wire \Selector3~1_combout ;
wire \Selector4~1_combout ;
wire \count[6]~15_combout ;
wire \count[0]~q ;
wire \count[0]~11 ;
wire \count[1]~12_combout ;
wire \count[1]~q ;
wire \count[1]~13 ;
wire \count[2]~16_combout ;
wire \count[2]~q ;
wire \count[2]~17 ;
wire \count[3]~18_combout ;
wire \count[3]~q ;
wire \max_reached~0_combout ;
wire \count[3]~19 ;
wire \count[4]~20_combout ;
wire \count[4]~q ;
wire \count[4]~21 ;
wire \count[5]~22_combout ;
wire \count[5]~q ;
wire \count[5]~23 ;
wire \count[6]~24_combout ;
wire \count[6]~q ;
wire \count[6]~25 ;
wire \count[7]~26_combout ;
wire \count[7]~q ;
wire \max_reached~1_combout ;
wire \count[7]~27 ;
wire \count[8]~28_combout ;
wire \count[8]~q ;
wire \count[8]~29 ;
wire \count[9]~30_combout ;
wire \count[9]~q ;
wire \max_reached~2_combout ;
wire \max_reached~3_combout ;
wire \max_reached~4_combout ;
wire \max_reached~q ;
wire \sink_comb_update_2~0_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~8_combout ;
wire \sink_state.run1~q ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \Selector5~2_combout ;
wire \sink_state.end1~q ;
wire \Selector0~0_combout ;
wire \sink_state.start~q ;
wire \Selector6~2_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;


fftsign_scfifo_1 \normal_fifo:fifo_eab_on:in_fifo (
	.q({q_unconnected_wire_21,q_unconnected_wire_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dffe_af(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.sink_out_stateempty_and_ready(\sink_out_state.empty_and_ready~q ),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(\sink_out_state.normal~q ),
	.sink_start(sink_start1),
	.empty_dff(empty_dff),
	.sink_stall(sink_stall1),
	.rdreq(\Selector7~0_combout ),
	.sink_staterun1(\sink_state.run1~q ),
	.sink_stateend1(\sink_state.end1~q ),
	.wrreq(\fifo_wrreq~0_combout ),
	.counter_reg_bit_0(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.data({gnd,gnd,\at_sink_data_int[19]~q ,\at_sink_data_int[18]~q ,\at_sink_data_int[17]~q ,\at_sink_data_int[16]~q ,\at_sink_data_int[15]~q ,\at_sink_data_int[14]~q ,\at_sink_data_int[13]~q ,\at_sink_data_int[12]~q ,\at_sink_data_int[11]~q ,\at_sink_data_int[10]~q ,
\at_sink_data_int[9]~q ,\at_sink_data_int[8]~q ,\at_sink_data_int[7]~q ,\at_sink_data_int[6]~q ,\at_sink_data_int[5]~q ,\at_sink_data_int[4]~q ,\at_sink_data_int[3]~q ,\at_sink_data_int[2]~q ,\at_sink_data_int[1]~q ,\at_sink_data_int[0]~q }),
	.clock(clk),
	.reset_n(reset_n));

cycloneive_lcell_comb \fifo_wrreq~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sink_state.run1~q ),
	.datad(\sink_state.end1~q ),
	.cin(gnd),
	.combout(\fifo_wrreq~0_combout ),
	.cout());
defparam \fifo_wrreq~0 .lut_mask = 16'h0FFF;
defparam \fifo_wrreq~0 .sum_lutc_input = "datac";

dffeas \at_sink_data_int[2] (
	.clk(clk),
	.d(at_sink_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[2]~q ),
	.prn(vcc));
defparam \at_sink_data_int[2] .is_wysiwyg = "true";
defparam \at_sink_data_int[2] .power_up = "low";

dffeas \at_sink_data_int[12] (
	.clk(clk),
	.d(at_sink_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[12]~q ),
	.prn(vcc));
defparam \at_sink_data_int[12] .is_wysiwyg = "true";
defparam \at_sink_data_int[12] .power_up = "low";

dffeas \at_sink_data_int[1] (
	.clk(clk),
	.d(at_sink_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[1]~q ),
	.prn(vcc));
defparam \at_sink_data_int[1] .is_wysiwyg = "true";
defparam \at_sink_data_int[1] .power_up = "low";

dffeas \at_sink_data_int[11] (
	.clk(clk),
	.d(at_sink_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[11]~q ),
	.prn(vcc));
defparam \at_sink_data_int[11] .is_wysiwyg = "true";
defparam \at_sink_data_int[11] .power_up = "low";

dffeas \at_sink_data_int[0] (
	.clk(clk),
	.d(at_sink_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[0]~q ),
	.prn(vcc));
defparam \at_sink_data_int[0] .is_wysiwyg = "true";
defparam \at_sink_data_int[0] .power_up = "low";

dffeas \at_sink_data_int[10] (
	.clk(clk),
	.d(at_sink_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[10]~q ),
	.prn(vcc));
defparam \at_sink_data_int[10] .is_wysiwyg = "true";
defparam \at_sink_data_int[10] .power_up = "low";

dffeas \at_sink_data_int[9] (
	.clk(clk),
	.d(at_sink_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[9]~q ),
	.prn(vcc));
defparam \at_sink_data_int[9] .is_wysiwyg = "true";
defparam \at_sink_data_int[9] .power_up = "low";

dffeas \at_sink_data_int[19] (
	.clk(clk),
	.d(at_sink_data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[19]~q ),
	.prn(vcc));
defparam \at_sink_data_int[19] .is_wysiwyg = "true";
defparam \at_sink_data_int[19] .power_up = "low";

dffeas \at_sink_data_int[8] (
	.clk(clk),
	.d(at_sink_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[8]~q ),
	.prn(vcc));
defparam \at_sink_data_int[8] .is_wysiwyg = "true";
defparam \at_sink_data_int[8] .power_up = "low";

dffeas \at_sink_data_int[18] (
	.clk(clk),
	.d(at_sink_data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[18]~q ),
	.prn(vcc));
defparam \at_sink_data_int[18] .is_wysiwyg = "true";
defparam \at_sink_data_int[18] .power_up = "low";

dffeas \at_sink_data_int[7] (
	.clk(clk),
	.d(at_sink_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[7]~q ),
	.prn(vcc));
defparam \at_sink_data_int[7] .is_wysiwyg = "true";
defparam \at_sink_data_int[7] .power_up = "low";

dffeas \at_sink_data_int[17] (
	.clk(clk),
	.d(at_sink_data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[17]~q ),
	.prn(vcc));
defparam \at_sink_data_int[17] .is_wysiwyg = "true";
defparam \at_sink_data_int[17] .power_up = "low";

dffeas \at_sink_data_int[6] (
	.clk(clk),
	.d(at_sink_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[6]~q ),
	.prn(vcc));
defparam \at_sink_data_int[6] .is_wysiwyg = "true";
defparam \at_sink_data_int[6] .power_up = "low";

dffeas \at_sink_data_int[16] (
	.clk(clk),
	.d(at_sink_data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[16]~q ),
	.prn(vcc));
defparam \at_sink_data_int[16] .is_wysiwyg = "true";
defparam \at_sink_data_int[16] .power_up = "low";

dffeas \at_sink_data_int[5] (
	.clk(clk),
	.d(at_sink_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[5]~q ),
	.prn(vcc));
defparam \at_sink_data_int[5] .is_wysiwyg = "true";
defparam \at_sink_data_int[5] .power_up = "low";

dffeas \at_sink_data_int[15] (
	.clk(clk),
	.d(at_sink_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[15]~q ),
	.prn(vcc));
defparam \at_sink_data_int[15] .is_wysiwyg = "true";
defparam \at_sink_data_int[15] .power_up = "low";

dffeas \at_sink_data_int[4] (
	.clk(clk),
	.d(at_sink_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[4]~q ),
	.prn(vcc));
defparam \at_sink_data_int[4] .is_wysiwyg = "true";
defparam \at_sink_data_int[4] .power_up = "low";

dffeas \at_sink_data_int[14] (
	.clk(clk),
	.d(at_sink_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[14]~q ),
	.prn(vcc));
defparam \at_sink_data_int[14] .is_wysiwyg = "true";
defparam \at_sink_data_int[14] .power_up = "low";

dffeas \at_sink_data_int[3] (
	.clk(clk),
	.d(at_sink_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[3]~q ),
	.prn(vcc));
defparam \at_sink_data_int[3] .is_wysiwyg = "true";
defparam \at_sink_data_int[3] .power_up = "low";

dffeas \at_sink_data_int[13] (
	.clk(clk),
	.d(at_sink_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[13]~q ),
	.prn(vcc));
defparam \at_sink_data_int[13] .is_wysiwyg = "true";
defparam \at_sink_data_int[13] .power_up = "low";

cycloneive_lcell_comb data_take(
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.end1~q ),
	.datac(\Selector2~8_combout ),
	.datad(\Selector4~1_combout ),
	.cin(gnd),
	.combout(\data_take~combout ),
	.cout());
defparam data_take.lut_mask = 16'hFFFE;
defparam data_take.sum_lutc_input = "datac";

dffeas at_sink_ready_s(
	.clk(clk),
	.d(\at_sink_ready_s~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_sink_ready_s1),
	.prn(vcc));
defparam at_sink_ready_s.is_wysiwyg = "true";
defparam at_sink_ready_s.power_up = "low";

dffeas send_eop_s(
	.clk(clk),
	.d(\Equal2~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_eop_s1),
	.prn(vcc));
defparam send_eop_s.is_wysiwyg = "true";
defparam send_eop_s.power_up = "low";

dffeas sink_start(
	.clk(clk),
	.d(\sink_start~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_start1),
	.prn(vcc));
defparam sink_start.is_wysiwyg = "true";
defparam sink_start.power_up = "low";

cycloneive_lcell_comb sink_stall(
	.dataa(gnd),
	.datab(gnd),
	.datac(sink_start1),
	.datad(empty_dff),
	.cin(gnd),
	.combout(sink_stall1),
	.cout());
defparam sink_stall.lut_mask = 16'h0FFF;
defparam sink_stall.sum_lutc_input = "datac";

dffeas \packet_error_s[1] (
	.clk(clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_1),
	.prn(vcc));
defparam \packet_error_s[1] .is_wysiwyg = "true";
defparam \packet_error_s[1] .power_up = "low";

dffeas \packet_error_s[0] (
	.clk(clk),
	.d(\Selector6~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_0),
	.prn(vcc));
defparam \packet_error_s[0] .is_wysiwyg = "true";
defparam \packet_error_s[0] .power_up = "low";

dffeas send_sop_s(
	.clk(clk),
	.d(\Equal1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_sop_s1),
	.prn(vcc));
defparam send_sop_s.is_wysiwyg = "true";
defparam send_sop_s.power_up = "low";

cycloneive_lcell_comb \at_sink_ready_s~0 (
	.dataa(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_sink_ready_s~0_combout ),
	.cout());
defparam \at_sink_ready_s~0 .lut_mask = 16'h5555;
defparam \at_sink_ready_s~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_cnt[0]~10 (
	.dataa(\out_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\out_cnt[0]~10_combout ),
	.cout(\out_cnt[0]~11 ));
defparam \out_cnt[0]~10 .lut_mask = 16'h55AA;
defparam \out_cnt[0]~10 .sum_lutc_input = "datac";

dffeas sink_stall_s(
	.clk(clk),
	.d(sink_stall1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_stall_s~q ),
	.prn(vcc));
defparam sink_stall_s.is_wysiwyg = "true";
defparam sink_stall_s.power_up = "low";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_stall_s~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFFF7;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \sink_out_state.normal (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.normal~q ),
	.prn(vcc));
defparam \sink_out_state.normal .is_wysiwyg = "true";
defparam \sink_out_state.normal .power_up = "low";

cycloneive_lcell_comb \Selector10~2 (
	.dataa(\sink_out_state.empty_and_ready~q ),
	.datab(sink_ready_ctrl),
	.datac(\sink_stall_s~q ),
	.datad(\sink_out_state.normal~q ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
defparam \Selector10~2 .lut_mask = 16'hBEFF;
defparam \Selector10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~3 (
	.dataa(sink_start1),
	.datab(empty_dff),
	.datac(\Selector10~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
defparam \Selector10~3 .lut_mask = 16'hF7F7;
defparam \Selector10~3 .sum_lutc_input = "datac";

dffeas \sink_out_state.empty_and_ready (
	.clk(clk),
	.d(\Selector10~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.empty_and_ready~q ),
	.prn(vcc));
defparam \sink_out_state.empty_and_ready .is_wysiwyg = "true";
defparam \sink_out_state.empty_and_ready .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\sink_out_state.empty_and_ready~q ),
	.datab(sink_ready_ctrl),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEFFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

cycloneive_lcell_comb \out_cnt[1]~12 (
	.dataa(\out_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[0]~11 ),
	.combout(\out_cnt[1]~12_combout ),
	.cout(\out_cnt[1]~13 ));
defparam \out_cnt[1]~12 .lut_mask = 16'h5A5F;
defparam \out_cnt[1]~12 .sum_lutc_input = "cin";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

cycloneive_lcell_comb \out_cnt[2]~14 (
	.dataa(\out_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[1]~13 ),
	.combout(\out_cnt[2]~14_combout ),
	.cout(\out_cnt[2]~15 ));
defparam \out_cnt[2]~14 .lut_mask = 16'h5AAF;
defparam \out_cnt[2]~14 .sum_lutc_input = "cin";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

cycloneive_lcell_comb \out_cnt[3]~16 (
	.dataa(\out_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[2]~15 ),
	.combout(\out_cnt[3]~16_combout ),
	.cout(\out_cnt[3]~17 ));
defparam \out_cnt[3]~16 .lut_mask = 16'h5A5F;
defparam \out_cnt[3]~16 .sum_lutc_input = "cin";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hFFFE;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_cnt[4]~18 (
	.dataa(\out_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[3]~17 ),
	.combout(\out_cnt[4]~18_combout ),
	.cout(\out_cnt[4]~19 ));
defparam \out_cnt[4]~18 .lut_mask = 16'h5AAF;
defparam \out_cnt[4]~18 .sum_lutc_input = "cin";

dffeas \out_cnt[4] (
	.clk(clk),
	.d(\out_cnt[4]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[4]~q ),
	.prn(vcc));
defparam \out_cnt[4] .is_wysiwyg = "true";
defparam \out_cnt[4] .power_up = "low";

cycloneive_lcell_comb \out_cnt[5]~20 (
	.dataa(\out_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[4]~19 ),
	.combout(\out_cnt[5]~20_combout ),
	.cout(\out_cnt[5]~21 ));
defparam \out_cnt[5]~20 .lut_mask = 16'h5A5F;
defparam \out_cnt[5]~20 .sum_lutc_input = "cin";

dffeas \out_cnt[5] (
	.clk(clk),
	.d(\out_cnt[5]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[5]~q ),
	.prn(vcc));
defparam \out_cnt[5] .is_wysiwyg = "true";
defparam \out_cnt[5] .power_up = "low";

cycloneive_lcell_comb \out_cnt[6]~22 (
	.dataa(\out_cnt[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[5]~21 ),
	.combout(\out_cnt[6]~22_combout ),
	.cout(\out_cnt[6]~23 ));
defparam \out_cnt[6]~22 .lut_mask = 16'h5AAF;
defparam \out_cnt[6]~22 .sum_lutc_input = "cin";

dffeas \out_cnt[6] (
	.clk(clk),
	.d(\out_cnt[6]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[6]~q ),
	.prn(vcc));
defparam \out_cnt[6] .is_wysiwyg = "true";
defparam \out_cnt[6] .power_up = "low";

cycloneive_lcell_comb \out_cnt[7]~24 (
	.dataa(\out_cnt[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[6]~23 ),
	.combout(\out_cnt[7]~24_combout ),
	.cout(\out_cnt[7]~25 ));
defparam \out_cnt[7]~24 .lut_mask = 16'h5A5F;
defparam \out_cnt[7]~24 .sum_lutc_input = "cin";

dffeas \out_cnt[7] (
	.clk(clk),
	.d(\out_cnt[7]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[7]~q ),
	.prn(vcc));
defparam \out_cnt[7] .is_wysiwyg = "true";
defparam \out_cnt[7] .power_up = "low";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hFFFE;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_cnt[8]~26 (
	.dataa(\out_cnt[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\out_cnt[7]~25 ),
	.combout(\out_cnt[8]~26_combout ),
	.cout(\out_cnt[8]~27 ));
defparam \out_cnt[8]~26 .lut_mask = 16'h5AAF;
defparam \out_cnt[8]~26 .sum_lutc_input = "cin";

dffeas \out_cnt[8] (
	.clk(clk),
	.d(\out_cnt[8]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[8]~q ),
	.prn(vcc));
defparam \out_cnt[8] .is_wysiwyg = "true";
defparam \out_cnt[8] .power_up = "low";

cycloneive_lcell_comb \out_cnt[9]~28 (
	.dataa(\out_cnt[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\out_cnt[8]~27 ),
	.combout(\out_cnt[9]~28_combout ),
	.cout());
defparam \out_cnt[9]~28 .lut_mask = 16'h5A5A;
defparam \out_cnt[9]~28 .sum_lutc_input = "cin";

dffeas \out_cnt[9] (
	.clk(clk),
	.d(\out_cnt[9]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\Equal2~2_combout ),
	.sload(gnd),
	.ena(\Selector7~0_combout ),
	.q(\out_cnt[9]~q ),
	.prn(vcc));
defparam \out_cnt[9] .is_wysiwyg = "true";
defparam \out_cnt[9] .power_up = "low";

cycloneive_lcell_comb \Equal2~2 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\out_cnt[8]~q ),
	.datad(\out_cnt[9]~q ),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hFFFE;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \send_sop_eop_p~0 (
	.dataa(sink_ready_ctrl),
	.datab(\sink_out_state.empty_and_ready~q ),
	.datac(\sink_out_state.normal~q ),
	.datad(sink_stall1),
	.cin(gnd),
	.combout(\send_sop_eop_p~0_combout ),
	.cout());
defparam \send_sop_eop_p~0 .lut_mask = 16'hEFFF;
defparam \send_sop_eop_p~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_start~0 (
	.dataa(sink_start1),
	.datab(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_start~0_combout ),
	.cout());
defparam \sink_start~0 .lut_mask = 16'hEEEE;
defparam \sink_start~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_comb_update_2~1 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sink_comb_update_2~1_combout ),
	.cout());
defparam \sink_comb_update_2~1 .lut_mask = 16'hEEEE;
defparam \sink_comb_update_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~10 (
	.dataa(\count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~10_combout ),
	.cout(\count[0]~11 ));
defparam \count[0]~10 .lut_mask = 16'h55AA;
defparam \count[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(at_sink_ready_s1),
	.datad(sink_valid),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hEFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \sink_state.stall (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.stall~q ),
	.prn(vcc));
defparam \sink_state.stall .is_wysiwyg = "true";
defparam \sink_state.stall .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sink_state.run1~q ),
	.datad(\sink_state.stall~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'h0FFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~6 (
	.dataa(sink_sop),
	.datab(\max_reached~q ),
	.datac(sink_eop),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hEFFF;
defparam \Selector2~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~7 (
	.dataa(sink_error_0),
	.datab(sink_error_1),
	.datac(\sink_comb_update_2~1_combout ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
defparam \Selector2~7 .lut_mask = 16'hFFFE;
defparam \Selector2~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_comb_update_2~2 (
	.dataa(at_sink_ready_s1),
	.datab(sink_eop),
	.datac(sink_valid),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~2_combout ),
	.cout());
defparam \sink_comb_update_2~2 .lut_mask = 16'hFEFF;
defparam \sink_comb_update_2~2 .sum_lutc_input = "datac";

dffeas \sink_state.st_err (
	.clk(clk),
	.d(\Selector3~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.st_err~q ),
	.prn(vcc));
defparam \sink_state.st_err .is_wysiwyg = "true";
defparam \sink_state.st_err .power_up = "low";

cycloneive_lcell_comb \Selector3~2 (
	.dataa(\sink_state.st_err~q ),
	.datab(\sink_comb_update_2~1_combout ),
	.datac(\Selector3~0_combout ),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hACFF;
defparam \Selector3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~2 (
	.dataa(\sink_comb_update_2~0_combout ),
	.datab(\sink_comb_update_2~1_combout ),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
defparam \Selector2~2 .lut_mask = 16'hFFFE;
defparam \Selector2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(sink_eop),
	.datab(sink_sop),
	.datac(sink_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'h7F7F;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~1 (
	.dataa(\max_reached~q ),
	.datab(sink_sop),
	.datac(at_sink_ready_s1),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hFFBF;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~3 (
	.dataa(\sink_state.run1~q ),
	.datab(at_sink_ready_s1),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
defparam \Selector2~3 .lut_mask = 16'hEDDE;
defparam \Selector2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~4 (
	.dataa(\sink_state.stall~q ),
	.datab(sink_valid),
	.datac(\sink_state.run1~q ),
	.datad(\Selector2~3_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
defparam \Selector2~4 .lut_mask = 16'hBFFB;
defparam \Selector2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~5 (
	.dataa(\Selector2~2_combout ),
	.datab(\Selector6~1_combout ),
	.datac(\Selector3~0_combout ),
	.datad(\Selector2~4_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
defparam \Selector2~5 .lut_mask = 16'hFFBF;
defparam \Selector2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~3 (
	.dataa(\Selector2~7_combout ),
	.datab(\sink_comb_update_2~2_combout ),
	.datac(\Selector3~2_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'hFAFC;
defparam \Selector3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[6]~14 (
	.dataa(\max_reached~q ),
	.datab(\Selector3~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[6]~14_combout ),
	.cout());
defparam \count[6]~14 .lut_mask = 16'hEEEE;
defparam \count[6]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(sink_error_0),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEFFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(gnd),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'hEEFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(sink_eop),
	.datab(\max_reached~q ),
	.datac(\Selector4~0_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFFFE;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[6]~15 (
	.dataa(\Selector2~8_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\Selector3~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[6]~15_combout ),
	.cout());
defparam \count[6]~15 .lut_mask = 16'hFEFE;
defparam \count[6]~15 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \count[1]~12 (
	.dataa(\count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~11 ),
	.combout(\count[1]~12_combout ),
	.cout(\count[1]~13 ));
defparam \count[1]~12 .lut_mask = 16'h5A5F;
defparam \count[1]~12 .sum_lutc_input = "cin";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \count[2]~16 (
	.dataa(\count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~13 ),
	.combout(\count[2]~16_combout ),
	.cout(\count[2]~17 ));
defparam \count[2]~16 .lut_mask = 16'h5AAF;
defparam \count[2]~16 .sum_lutc_input = "cin";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count[3]~18 (
	.dataa(\count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~17 ),
	.combout(\count[3]~18_combout ),
	.cout(\count[3]~19 ));
defparam \count[3]~18 .lut_mask = 16'h5A5F;
defparam \count[3]~18 .sum_lutc_input = "cin";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \max_reached~0 (
	.dataa(\count[1]~q ),
	.datab(\count[2]~q ),
	.datac(\count[3]~q ),
	.datad(\count[0]~q ),
	.cin(gnd),
	.combout(\max_reached~0_combout ),
	.cout());
defparam \max_reached~0 .lut_mask = 16'hFEFF;
defparam \max_reached~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[4]~20 (
	.dataa(\count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~19 ),
	.combout(\count[4]~20_combout ),
	.cout(\count[4]~21 ));
defparam \count[4]~20 .lut_mask = 16'h5AAF;
defparam \count[4]~20 .sum_lutc_input = "cin";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count[5]~22 (
	.dataa(\count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~21 ),
	.combout(\count[5]~22_combout ),
	.cout(\count[5]~23 ));
defparam \count[5]~22 .lut_mask = 16'h5A5F;
defparam \count[5]~22 .sum_lutc_input = "cin";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count[6]~24 (
	.dataa(\count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~23 ),
	.combout(\count[6]~24_combout ),
	.cout(\count[6]~25 ));
defparam \count[6]~24 .lut_mask = 16'h5AAF;
defparam \count[6]~24 .sum_lutc_input = "cin";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count[7]~26 (
	.dataa(\count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~25 ),
	.combout(\count[7]~26_combout ),
	.cout(\count[7]~27 ));
defparam \count[7]~26 .lut_mask = 16'h5A5F;
defparam \count[7]~26 .sum_lutc_input = "cin";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \max_reached~1 (
	.dataa(\count[4]~q ),
	.datab(\count[5]~q ),
	.datac(\count[6]~q ),
	.datad(\count[7]~q ),
	.cin(gnd),
	.combout(\max_reached~1_combout ),
	.cout());
defparam \max_reached~1 .lut_mask = 16'hFFFE;
defparam \max_reached~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[8]~28 (
	.dataa(\count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[7]~27 ),
	.combout(\count[8]~28_combout ),
	.cout(\count[8]~29 ));
defparam \count[8]~28 .lut_mask = 16'h5AAF;
defparam \count[8]~28 .sum_lutc_input = "cin";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \count[9]~30 (
	.dataa(\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[8]~29 ),
	.combout(\count[9]~30_combout ),
	.cout());
defparam \count[9]~30 .lut_mask = 16'h5A5A;
defparam \count[9]~30 .sum_lutc_input = "cin";

dffeas \count[9] (
	.clk(clk),
	.d(\count[9]~30_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\count[6]~14_combout ),
	.sload(gnd),
	.ena(\count[6]~15_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \max_reached~2 (
	.dataa(\max_reached~0_combout ),
	.datab(\max_reached~1_combout ),
	.datac(\count[8]~q ),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\max_reached~2_combout ),
	.cout());
defparam \max_reached~2 .lut_mask = 16'hFFFE;
defparam \max_reached~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \max_reached~3 (
	.dataa(\Selector2~8_combout ),
	.datab(\Selector4~1_combout ),
	.datac(gnd),
	.datad(\Selector3~3_combout ),
	.cin(gnd),
	.combout(\max_reached~3_combout ),
	.cout());
defparam \max_reached~3 .lut_mask = 16'hEEFF;
defparam \max_reached~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \max_reached~4 (
	.dataa(\max_reached~2_combout ),
	.datab(\max_reached~q ),
	.datac(gnd),
	.datad(\max_reached~3_combout ),
	.cin(gnd),
	.combout(\max_reached~4_combout ),
	.cout());
defparam \max_reached~4 .lut_mask = 16'hAACC;
defparam \max_reached~4 .sum_lutc_input = "datac";

dffeas max_reached(
	.clk(clk),
	.d(\max_reached~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\max_reached~q ),
	.prn(vcc));
defparam max_reached.is_wysiwyg = "true";
defparam max_reached.power_up = "low";

cycloneive_lcell_comb \sink_comb_update_2~0 (
	.dataa(at_sink_ready_s1),
	.datab(sink_valid),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\sink_comb_update_2~0_combout ),
	.cout());
defparam \sink_comb_update_2~0 .lut_mask = 16'hEFFF;
defparam \sink_comb_update_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(sink_sop),
	.datab(sink_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEEEE;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~1 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(at_sink_ready_s1),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFFFB;
defparam \Selector2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~8 (
	.dataa(\sink_comb_update_2~0_combout ),
	.datab(\Selector2~1_combout ),
	.datac(\Selector2~5_combout ),
	.datad(\Selector2~7_combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
defparam \Selector2~8 .lut_mask = 16'hACFF;
defparam \Selector2~8 .sum_lutc_input = "datac";

dffeas \sink_state.run1 (
	.clk(clk),
	.d(\Selector2~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.run1~q ),
	.prn(vcc));
defparam \sink_state.run1 .is_wysiwyg = "true";
defparam \sink_state.run1 .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\sink_state.run1~q ),
	.datab(\sink_state.stall~q ),
	.datac(sink_eop),
	.datad(\max_reached~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEFFE;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(sink_sop),
	.datad(sink_error_0),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'h0FFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~2 (
	.dataa(\sink_comb_update_2~1_combout ),
	.datab(sink_error_1),
	.datac(\Selector5~0_combout ),
	.datad(\Selector5~1_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hFFFE;
defparam \Selector5~2 .sum_lutc_input = "datac";

dffeas \sink_state.end1 (
	.clk(clk),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.end1~q ),
	.prn(vcc));
defparam \sink_state.end1 .is_wysiwyg = "true";
defparam \sink_state.end1 .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\sink_state.end1~q ),
	.datab(\sink_state.st_err~q ),
	.datac(\sink_state.start~q ),
	.datad(\sink_comb_update_2~1_combout ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFFF7;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \sink_state.start (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.start~q ),
	.prn(vcc));
defparam \sink_state.start .is_wysiwyg = "true";
defparam \sink_state.start .power_up = "low";

cycloneive_lcell_comb \Selector6~2 (
	.dataa(\sink_state.end1~q ),
	.datab(\sink_state.st_err~q ),
	.datac(gnd),
	.datad(\sink_state.start~q ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hEEFF;
defparam \Selector6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~3 (
	.dataa(\Selector3~1_combout ),
	.datab(\Selector6~2_combout ),
	.datac(\Selector3~0_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
defparam \Selector6~3 .lut_mask = 16'hEFFF;
defparam \Selector6~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~4 (
	.dataa(sink_error_0),
	.datab(\Selector6~3_combout ),
	.datac(\sink_comb_update_2~1_combout ),
	.datad(sink_error_1),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
defparam \Selector6~4 .lut_mask = 16'hACFF;
defparam \Selector6~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h7FFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(\out_cnt[4]~q ),
	.datab(\out_cnt[5]~q ),
	.datac(\out_cnt[6]~q ),
	.datad(\out_cnt[7]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h7FFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\out_cnt[8]~q ),
	.datad(\out_cnt[9]~q ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hEFFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

endmodule

module fftsign_scfifo_1 (
	q,
	dffe_af,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff,
	sink_stall,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
output 	dffe_af;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff;
input 	sink_stall;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[21:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fftsign_scfifo_o2j1 auto_generated(
	.q({q_unconnected_wire_21,q_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.dffe_af1(dffe_af),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(sink_out_statenormal),
	.sink_start(sink_start),
	.empty_dff(empty_dff),
	.sink_stall(sink_stall),
	.rdreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wrreq(wrreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	.data({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module fftsign_scfifo_o2j1 (
	q,
	dffe_af1,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff,
	sink_stall,
	rdreq,
	sink_staterun1,
	sink_stateend1,
	wrreq,
	counter_reg_bit_0,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
output 	dffe_af1;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff;
input 	sink_stall;
input 	rdreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wrreq;
output 	counter_reg_bit_0;
input 	[21:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;


fftsign_a_dpfifo_cc81 dpfifo(
	.q({q_unconnected_wire_21,q_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_out_statenormal(sink_out_statenormal),
	.sink_start(sink_start),
	.empty_dff1(empty_dff),
	.sink_stall(sink_stall),
	.rreq(rdreq),
	.sink_staterun1(sink_staterun1),
	.sink_stateend1(sink_stateend1),
	.wreq(wrreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	.data({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock),
	.reset_n(reset_n));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

cycloneive_lcell_comb \dffe_af~0 (
	.dataa(rdreq),
	.datab(wrreq),
	.datac(dffe_af1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\dffe_af~0_combout ),
	.cout());
defparam \dffe_af~0 .lut_mask = 16'hF7FF;
defparam \dffe_af~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_af~1 (
	.dataa(dffe_af1),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datad(\dffe_af~0_combout ),
	.cin(gnd),
	.combout(\dffe_af~1_combout ),
	.cout());
defparam \dffe_af~1 .lut_mask = 16'hFFBE;
defparam \dffe_af~1 .sum_lutc_input = "datac";

endmodule

module fftsign_a_dpfifo_cc81 (
	q,
	counter_reg_bit_2,
	counter_reg_bit_1,
	sink_out_stateempty_and_ready,
	sink_ready_ctrl,
	sink_out_statenormal,
	sink_start,
	empty_dff1,
	sink_stall,
	rreq,
	sink_staterun1,
	sink_stateend1,
	wreq,
	counter_reg_bit_0,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	sink_out_stateempty_and_ready;
input 	sink_ready_ctrl;
input 	sink_out_statenormal;
input 	sink_start;
output 	empty_dff1;
input 	sink_stall;
input 	rreq;
input 	sink_staterun1;
input 	sink_stateend1;
input 	wreq;
output 	counter_reg_bit_0;
input 	[21:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \_~8_combout ;
wire \_~9_combout ;
wire \_~10_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \_~5_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_is_1_dff~q ;
wire \_~7_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_will_be_1~0_combout ;
wire \_~6_combout ;
wire \_~11_combout ;


fftsign_cntr_unb wr_ptr(
	.fifo_wrreq(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.clock(clock),
	.reset_n(reset_n));

fftsign_cntr_ao7 usedw_counter(
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.updown(wreq),
	.counter_reg_bit_0(counter_reg_bit_0),
	._(\_~4_combout ),
	.clock(clock),
	.reset_n(reset_n));

fftsign_cntr_tnb rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	._(\_~9_combout ),
	.clock(clock),
	.reset_n(reset_n));

fftsign_altsyncram_g8j1 FIFOram(
	.q_b({q_b_unconnected_wire_21,q_b_unconnected_wire_20,q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(rreq),
	.wren_a(wreq),
	.data_a({gnd,gnd,data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

cycloneive_lcell_comb \_~4 (
	.dataa(wreq),
	.datab(sink_out_stateempty_and_ready),
	.datac(sink_ready_ctrl),
	.datad(\_~10_combout ),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h6996;
defparam \_~4 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rreq),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(rreq),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(rreq),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~8 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(sink_out_stateempty_and_ready),
	.datac(sink_out_statenormal),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~8_combout ),
	.cout());
defparam \_~8 .lut_mask = 16'hDFDF;
defparam \_~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~9 (
	.dataa(sink_out_stateempty_and_ready),
	.datab(sink_ready_ctrl),
	.datac(sink_stall),
	.datad(\_~8_combout ),
	.cin(gnd),
	.combout(\_~9_combout ),
	.cout());
defparam \_~9 .lut_mask = 16'hFFEF;
defparam \_~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~10 (
	.dataa(sink_start),
	.datab(empty_dff1),
	.datac(sink_out_stateempty_and_ready),
	.datad(sink_out_statenormal),
	.cin(gnd),
	.combout(\_~10_combout ),
	.cout());
defparam \_~10 .lut_mask = 16'hFEFF;
defparam \_~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'h5555;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\_~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \_~5 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(counter_reg_bit_0),
	.datad(counter_reg_bit_2),
	.cin(gnd),
	.combout(\_~5_combout ),
	.cout());
defparam \_~5 .lut_mask = 16'hAFFF;
defparam \_~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_will_be_1~0_combout ),
	.datab(\usedw_is_1_dff~q ),
	.datac(rreq),
	.datad(wreq),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hEFFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \_~7 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(rreq),
	.datac(wreq),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\_~7_combout ),
	.cout());
defparam \_~7 .lut_mask = 16'hFF7D;
defparam \_~7 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\_~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~5_combout ),
	.datab(rreq),
	.datac(wreq),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBEFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~6 (
	.dataa(wreq),
	.datab(\usedw_is_1_dff~q ),
	.datac(rreq),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\_~6_combout ),
	.cout());
defparam \_~6 .lut_mask = 16'hDEFF;
defparam \_~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~11 (
	.dataa(sink_staterun1),
	.datab(sink_stateend1),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\_~6_combout ),
	.cin(gnd),
	.combout(\_~11_combout ),
	.cout());
defparam \_~11 .lut_mask = 16'h7FFF;
defparam \_~11 .sum_lutc_input = "datac";

endmodule

module fftsign_altsyncram_g8j1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[21:0] data_a;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 22;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 22;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 22;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 22;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 22;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 22;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 3;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 7;
defparam ram_block1a19.port_a_logical_ram_depth = 8;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 3;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 7;
defparam ram_block1a18.port_a_logical_ram_depth = 8;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 3;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 7;
defparam ram_block1a17.port_a_logical_ram_depth = 8;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 3;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 7;
defparam ram_block1a16.port_a_logical_ram_depth = 8;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 22;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 22;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 22;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 22;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "fftsign_fft_ii_0:fft_ii_0|asj_fft_si_se_so_b:asj_fft_si_se_so_b_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_o2j1:auto_generated|a_dpfifo_cc81:dpfifo|altsyncram_g8j1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

endmodule

module fftsign_cntr_ao7 (
	counter_reg_bit_2,
	counter_reg_bit_1,
	updown,
	counter_reg_bit_0,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	updown;
output 	counter_reg_bit_0;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fftsign_cntr_tnb (
	counter_reg_bit_0,
	counter_reg_bit_1,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout());
defparam counter_comb_bita1.lut_mask = 16'h5A5A;
defparam counter_comb_bita1.sum_lutc_input = "cin";

endmodule

module fftsign_cntr_unb (
	fifo_wrreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	fifo_wrreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module fftsign_auk_dspip_avalon_streaming_source (
	data_count,
	at_source_valid_s1,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s1,
	at_source_eop_s1,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_22,
	at_source_data_23,
	at_source_data_24,
	at_source_data_25,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_14,
	at_source_data_15,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	source_packet_error_1,
	source_packet_error_0,
	source_stall_reg,
	sink_stall_reg,
	master_source_ena,
	sink_ready_ctrl_d,
	send_sop_s,
	sop,
	global_clock_enable,
	stall_reg,
	source_stall_int_d1,
	data,
	Mux0,
	clk,
	reset_n,
	source_ready)/* synthesis synthesis_greybox=1 */;
input 	[9:0] data_count;
output 	at_source_valid_s1;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s1;
output 	at_source_eop_s1;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_22;
output 	at_source_data_23;
output 	at_source_data_24;
output 	at_source_data_25;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
input 	source_packet_error_1;
input 	source_packet_error_0;
input 	source_stall_reg;
input 	sink_stall_reg;
input 	master_source_ena;
input 	sink_ready_ctrl_d;
input 	send_sop_s;
input 	sop;
input 	global_clock_enable;
input 	stall_reg;
output 	source_stall_int_d1;
input 	[25:0] data;
output 	Mux0;
input 	clk;
input 	reset_n;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_multi:source_state.end1~q ;
wire \packet_error0~combout ;
wire \Selector3~0_combout ;
wire \stall_controller_comb~0_combout ;
wire \was_stalled~1_combout ;
wire \was_stalled~0_combout ;
wire \was_stalled~2_combout ;
wire \was_stalled~q ;
wire \stall_controller_comb~1_combout ;
wire \Mux1~0_combout ;
wire \valid_ctrl_inter~0_combout ;
wire \data_wr_enb0~0_combout ;
wire \Mux2~1_combout ;
wire \valid_ctrl_inter~1_combout ;
wire \valid_ctrl_int~q ;
wire \Mux2~0_combout ;
wire \Mux3~0_combout ;
wire \valid_ctrl_inter1~0_combout ;
wire \valid_ctrl_int1~q ;
wire \first_data~0_combout ;
wire \first_data~q ;
wire \data_select~0_combout ;
wire \data_count_int1[7]~q ;
wire \data_count_int[9]~q ;
wire \data_count_int[7]~q ;
wire \data_count_int[8]~q ;
wire \data_count_int[3]~q ;
wire \packet_multi:count_finished~0_combout ;
wire \data_count_int1[9]~q ;
wire \data_count_int1[8]~q ;
wire \data_count_int1[3]~q ;
wire \packet_multi:count_finished~1_combout ;
wire \packet_multi:count_finished~2_combout ;
wire \data_count_int1[4]~q ;
wire \data_count_int[4]~q ;
wire \data_count_int[6]~q ;
wire \data_count_int[5]~q ;
wire \data_count_int[2]~q ;
wire \packet_multi:count_finished~3_combout ;
wire \data_count_int1[6]~q ;
wire \data_count_int1[5]~q ;
wire \data_count_int1[2]~q ;
wire \packet_multi:count_finished~4_combout ;
wire \packet_multi:count_finished~5_combout ;
wire \data_count_int[0]~q ;
wire \data_count_int1[0]~q ;
wire \data_count_int1[1]~q ;
wire \data_count_int[1]~q ;
wire \data_count_int_selected[1]~0_combout ;
wire \packet_multi:count_finished~6_combout ;
wire \at_source_valid_int~0_combout ;
wire \packet_multi:count_finished~combout ;
wire \Selector1~1_combout ;
wire \Selector1~0_combout ;
wire \Selector1~2_combout ;
wire \source_comb_update_2~0_combout ;
wire \source_comb_update_2~1_combout ;
wire \source_comb_update_2~2_combout ;
wire \source_comb_update_2~3_combout ;
wire \source_comb_update_2~4_combout ;
wire \source_comb_update_2~5_combout ;
wire \source_comb_update_2~6_combout ;
wire \source_comb_update_2~7_combout ;
wire \Selector1~3_combout ;
wire \packet_multi:source_state.st_err~q ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \packet_multi:source_state.start~q ;
wire \Selector1~4_combout ;
wire \Selector1~5_combout ;
wire \packet_multi:source_state.sop~q ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \packet_multi:source_state.run1~q ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \at_source_valid_int~1_combout ;
wire \at_source_valid_int~2_combout ;
wire \at_source_valid_int~3_combout ;
wire \at_source_valid_int~4_combout ;
wire \Selector5~0_combout ;
wire \Selector2~6_combout ;
wire \Selector5~1_combout ;
wire \data_int1[16]~q ;
wire \data_int[16]~q ;
wire \data_int_selected[16]~0_combout ;
wire \data_int1[17]~q ;
wire \data_int[17]~q ;
wire \data_int_selected[17]~1_combout ;
wire \data_int1[18]~q ;
wire \data_int[18]~q ;
wire \data_int_selected[18]~2_combout ;
wire \data_int1[19]~q ;
wire \data_int[19]~q ;
wire \data_int_selected[19]~3_combout ;
wire \data_int1[20]~q ;
wire \data_int[20]~q ;
wire \data_int_selected[20]~4_combout ;
wire \data_int1[21]~q ;
wire \data_int[21]~q ;
wire \data_int_selected[21]~5_combout ;
wire \data_int1[22]~q ;
wire \data_int[22]~q ;
wire \data_int_selected[22]~6_combout ;
wire \data_int1[23]~q ;
wire \data_int[23]~q ;
wire \data_int_selected[23]~7_combout ;
wire \data_int1[24]~q ;
wire \data_int[24]~q ;
wire \data_int_selected[24]~8_combout ;
wire \data_int1[25]~q ;
wire \data_int[25]~q ;
wire \data_int_selected[25]~9_combout ;
wire \data_int1[6]~q ;
wire \data_int[6]~q ;
wire \data_int_selected[6]~10_combout ;
wire \data_int1[7]~q ;
wire \data_int[7]~q ;
wire \data_int_selected[7]~11_combout ;
wire \data_int1[8]~q ;
wire \data_int[8]~q ;
wire \data_int_selected[8]~12_combout ;
wire \data_int1[9]~q ;
wire \data_int[9]~q ;
wire \data_int_selected[9]~13_combout ;
wire \data_int1[10]~q ;
wire \data_int[10]~q ;
wire \data_int_selected[10]~14_combout ;
wire \data_int1[11]~q ;
wire \data_int[11]~q ;
wire \data_int_selected[11]~15_combout ;
wire \data_int1[12]~q ;
wire \data_int[12]~q ;
wire \data_int_selected[12]~16_combout ;
wire \data_int1[13]~q ;
wire \data_int[13]~q ;
wire \data_int_selected[13]~17_combout ;
wire \data_int1[14]~q ;
wire \data_int[14]~q ;
wire \data_int_selected[14]~18_combout ;
wire \data_int1[15]~q ;
wire \data_int[15]~q ;
wire \data_int_selected[15]~19_combout ;
wire \data_int1[0]~q ;
wire \data_int[0]~q ;
wire \data_int_selected[0]~20_combout ;
wire \data_int1[1]~q ;
wire \data_int[1]~q ;
wire \data_int_selected[1]~21_combout ;
wire \data_int1[2]~q ;
wire \data_int[2]~q ;
wire \data_int_selected[2]~22_combout ;
wire \data_int1[3]~q ;
wire \data_int[3]~q ;
wire \data_int_selected[3]~23_combout ;
wire \data_int1[4]~q ;
wire \data_int[4]~q ;
wire \data_int_selected[4]~24_combout ;
wire \data_int1[5]~q ;
wire \data_int[5]~q ;
wire \data_int_selected[5]~25_combout ;
wire \Mux0~0_combout ;


dffeas at_source_valid_s(
	.clk(clk),
	.d(\at_source_valid_int~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_valid_s1),
	.prn(vcc));
defparam at_source_valid_s.is_wysiwyg = "true";
defparam at_source_valid_s.power_up = "low";

dffeas \at_source_error[0] (
	.clk(clk),
	.d(source_packet_error_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_0),
	.prn(vcc));
defparam \at_source_error[0] .is_wysiwyg = "true";
defparam \at_source_error[0] .power_up = "low";

dffeas \at_source_error[1] (
	.clk(clk),
	.d(source_packet_error_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_1),
	.prn(vcc));
defparam \at_source_error[1] .is_wysiwyg = "true";
defparam \at_source_error[1] .power_up = "low";

dffeas at_source_sop_s(
	.clk(clk),
	.d(\Selector1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_sop_s1),
	.prn(vcc));
defparam at_source_sop_s.is_wysiwyg = "true";
defparam at_source_sop_s.power_up = "low";

dffeas at_source_eop_s(
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_eop_s1),
	.prn(vcc));
defparam at_source_eop_s.is_wysiwyg = "true";
defparam at_source_eop_s.power_up = "low";

dffeas \at_source_data[16] (
	.clk(clk),
	.d(\data_int_selected[16]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_16),
	.prn(vcc));
defparam \at_source_data[16] .is_wysiwyg = "true";
defparam \at_source_data[16] .power_up = "low";

dffeas \at_source_data[17] (
	.clk(clk),
	.d(\data_int_selected[17]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_17),
	.prn(vcc));
defparam \at_source_data[17] .is_wysiwyg = "true";
defparam \at_source_data[17] .power_up = "low";

dffeas \at_source_data[18] (
	.clk(clk),
	.d(\data_int_selected[18]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_18),
	.prn(vcc));
defparam \at_source_data[18] .is_wysiwyg = "true";
defparam \at_source_data[18] .power_up = "low";

dffeas \at_source_data[19] (
	.clk(clk),
	.d(\data_int_selected[19]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_19),
	.prn(vcc));
defparam \at_source_data[19] .is_wysiwyg = "true";
defparam \at_source_data[19] .power_up = "low";

dffeas \at_source_data[20] (
	.clk(clk),
	.d(\data_int_selected[20]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_20),
	.prn(vcc));
defparam \at_source_data[20] .is_wysiwyg = "true";
defparam \at_source_data[20] .power_up = "low";

dffeas \at_source_data[21] (
	.clk(clk),
	.d(\data_int_selected[21]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_21),
	.prn(vcc));
defparam \at_source_data[21] .is_wysiwyg = "true";
defparam \at_source_data[21] .power_up = "low";

dffeas \at_source_data[22] (
	.clk(clk),
	.d(\data_int_selected[22]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_22),
	.prn(vcc));
defparam \at_source_data[22] .is_wysiwyg = "true";
defparam \at_source_data[22] .power_up = "low";

dffeas \at_source_data[23] (
	.clk(clk),
	.d(\data_int_selected[23]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_23),
	.prn(vcc));
defparam \at_source_data[23] .is_wysiwyg = "true";
defparam \at_source_data[23] .power_up = "low";

dffeas \at_source_data[24] (
	.clk(clk),
	.d(\data_int_selected[24]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_24),
	.prn(vcc));
defparam \at_source_data[24] .is_wysiwyg = "true";
defparam \at_source_data[24] .power_up = "low";

dffeas \at_source_data[25] (
	.clk(clk),
	.d(\data_int_selected[25]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_25),
	.prn(vcc));
defparam \at_source_data[25] .is_wysiwyg = "true";
defparam \at_source_data[25] .power_up = "low";

dffeas \at_source_data[6] (
	.clk(clk),
	.d(\data_int_selected[6]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_6),
	.prn(vcc));
defparam \at_source_data[6] .is_wysiwyg = "true";
defparam \at_source_data[6] .power_up = "low";

dffeas \at_source_data[7] (
	.clk(clk),
	.d(\data_int_selected[7]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_7),
	.prn(vcc));
defparam \at_source_data[7] .is_wysiwyg = "true";
defparam \at_source_data[7] .power_up = "low";

dffeas \at_source_data[8] (
	.clk(clk),
	.d(\data_int_selected[8]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_8),
	.prn(vcc));
defparam \at_source_data[8] .is_wysiwyg = "true";
defparam \at_source_data[8] .power_up = "low";

dffeas \at_source_data[9] (
	.clk(clk),
	.d(\data_int_selected[9]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_9),
	.prn(vcc));
defparam \at_source_data[9] .is_wysiwyg = "true";
defparam \at_source_data[9] .power_up = "low";

dffeas \at_source_data[10] (
	.clk(clk),
	.d(\data_int_selected[10]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_10),
	.prn(vcc));
defparam \at_source_data[10] .is_wysiwyg = "true";
defparam \at_source_data[10] .power_up = "low";

dffeas \at_source_data[11] (
	.clk(clk),
	.d(\data_int_selected[11]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_11),
	.prn(vcc));
defparam \at_source_data[11] .is_wysiwyg = "true";
defparam \at_source_data[11] .power_up = "low";

dffeas \at_source_data[12] (
	.clk(clk),
	.d(\data_int_selected[12]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_12),
	.prn(vcc));
defparam \at_source_data[12] .is_wysiwyg = "true";
defparam \at_source_data[12] .power_up = "low";

dffeas \at_source_data[13] (
	.clk(clk),
	.d(\data_int_selected[13]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_13),
	.prn(vcc));
defparam \at_source_data[13] .is_wysiwyg = "true";
defparam \at_source_data[13] .power_up = "low";

dffeas \at_source_data[14] (
	.clk(clk),
	.d(\data_int_selected[14]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_14),
	.prn(vcc));
defparam \at_source_data[14] .is_wysiwyg = "true";
defparam \at_source_data[14] .power_up = "low";

dffeas \at_source_data[15] (
	.clk(clk),
	.d(\data_int_selected[15]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_15),
	.prn(vcc));
defparam \at_source_data[15] .is_wysiwyg = "true";
defparam \at_source_data[15] .power_up = "low";

dffeas \at_source_data[0] (
	.clk(clk),
	.d(\data_int_selected[0]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_0),
	.prn(vcc));
defparam \at_source_data[0] .is_wysiwyg = "true";
defparam \at_source_data[0] .power_up = "low";

dffeas \at_source_data[1] (
	.clk(clk),
	.d(\data_int_selected[1]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_1),
	.prn(vcc));
defparam \at_source_data[1] .is_wysiwyg = "true";
defparam \at_source_data[1] .power_up = "low";

dffeas \at_source_data[2] (
	.clk(clk),
	.d(\data_int_selected[2]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_2),
	.prn(vcc));
defparam \at_source_data[2] .is_wysiwyg = "true";
defparam \at_source_data[2] .power_up = "low";

dffeas \at_source_data[3] (
	.clk(clk),
	.d(\data_int_selected[3]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_3),
	.prn(vcc));
defparam \at_source_data[3] .is_wysiwyg = "true";
defparam \at_source_data[3] .power_up = "low";

dffeas \at_source_data[4] (
	.clk(clk),
	.d(\data_int_selected[4]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_4),
	.prn(vcc));
defparam \at_source_data[4] .is_wysiwyg = "true";
defparam \at_source_data[4] .power_up = "low";

dffeas \at_source_data[5] (
	.clk(clk),
	.d(\data_int_selected[5]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_5),
	.prn(vcc));
defparam \at_source_data[5] .is_wysiwyg = "true";
defparam \at_source_data[5] .power_up = "low";

dffeas source_stall_int_d(
	.clk(clk),
	.d(Mux0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_int_d1),
	.prn(vcc));
defparam source_stall_int_d.is_wysiwyg = "true";
defparam source_stall_int_d.power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\valid_ctrl_int~q ),
	.datab(\stall_controller_comb~1_combout ),
	.datac(\valid_ctrl_int1~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFFE;
defparam \Mux0~1 .sum_lutc_input = "datac";

dffeas \packet_multi:source_state.end1 (
	.clk(clk),
	.d(\Selector3~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.end1~q ),
	.prn(vcc));
defparam \packet_multi:source_state.end1 .is_wysiwyg = "true";
defparam \packet_multi:source_state.end1 .power_up = "low";

cycloneive_lcell_comb packet_error0(
	.dataa(source_packet_error_1),
	.datab(source_packet_error_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_error0~combout ),
	.cout());
defparam packet_error0.lut_mask = 16'hEEEE;
defparam packet_error0.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\packet_multi:source_state.end1~q ),
	.datab(at_source_valid_s1),
	.datac(source_ready),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hBFFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \stall_controller_comb~0 (
	.dataa(sink_stall_reg),
	.datab(sink_ready_ctrl_d),
	.datac(send_sop_s),
	.datad(sop),
	.cin(gnd),
	.combout(\stall_controller_comb~0_combout ),
	.cout());
defparam \stall_controller_comb~0 .lut_mask = 16'hBFFF;
defparam \stall_controller_comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \was_stalled~1 (
	.dataa(source_ready),
	.datab(\first_data~q ),
	.datac(at_source_valid_s1),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\was_stalled~1_combout ),
	.cout());
defparam \was_stalled~1 .lut_mask = 16'hEFFF;
defparam \was_stalled~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \was_stalled~0 (
	.dataa(global_clock_enable),
	.datab(stall_reg),
	.datac(gnd),
	.datad(source_stall_int_d1),
	.cin(gnd),
	.combout(\was_stalled~0_combout ),
	.cout());
defparam \was_stalled~0 .lut_mask = 16'hEEFF;
defparam \was_stalled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \was_stalled~2 (
	.dataa(\was_stalled~q ),
	.datab(\stall_controller_comb~1_combout ),
	.datac(\was_stalled~1_combout ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\was_stalled~2_combout ),
	.cout());
defparam \was_stalled~2 .lut_mask = 16'hFEFF;
defparam \was_stalled~2 .sum_lutc_input = "datac";

dffeas was_stalled(
	.clk(clk),
	.d(\was_stalled~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\was_stalled~q ),
	.prn(vcc));
defparam was_stalled.is_wysiwyg = "true";
defparam was_stalled.power_up = "low";

cycloneive_lcell_comb \stall_controller_comb~1 (
	.dataa(master_source_ena),
	.datab(\stall_controller_comb~0_combout ),
	.datac(source_stall_reg),
	.datad(\was_stalled~q ),
	.cin(gnd),
	.combout(\stall_controller_comb~1_combout ),
	.cout());
defparam \stall_controller_comb~1 .lut_mask = 16'hEFFF;
defparam \stall_controller_comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(source_ready),
	.datab(\valid_ctrl_int1~q ),
	.datac(\valid_ctrl_int~q ),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFAFC;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_inter~0 (
	.dataa(\valid_ctrl_int~q ),
	.datab(\data_select~0_combout ),
	.datac(\Mux1~0_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~0_combout ),
	.cout());
defparam \valid_ctrl_inter~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_wr_enb0~0 (
	.dataa(source_ready),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\data_wr_enb0~0_combout ),
	.cout());
defparam \data_wr_enb0~0 .lut_mask = 16'hFEFF;
defparam \data_wr_enb0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\stall_controller_comb~1_combout ),
	.datab(\data_wr_enb0~0_combout ),
	.datac(gnd),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hEEFF;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_inter~1 (
	.dataa(\valid_ctrl_inter~0_combout ),
	.datab(\Mux2~1_combout ),
	.datac(\was_stalled~q ),
	.datad(\was_stalled~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter~1_combout ),
	.cout());
defparam \valid_ctrl_inter~1 .lut_mask = 16'h8BFF;
defparam \valid_ctrl_inter~1 .sum_lutc_input = "datac";

dffeas valid_ctrl_int(
	.clk(clk),
	.d(\valid_ctrl_inter~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int~q ),
	.prn(vcc));
defparam valid_ctrl_int.is_wysiwyg = "true";
defparam valid_ctrl_int.power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(at_source_valid_s1),
	.datab(\valid_ctrl_int1~q ),
	.datac(\valid_ctrl_int~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFEFE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\stall_controller_comb~1_combout ),
	.datab(\Mux2~0_combout ),
	.datac(source_ready),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hEFFF;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_ctrl_inter1~0 (
	.dataa(\Mux3~0_combout ),
	.datab(\valid_ctrl_int1~q ),
	.datac(\data_select~0_combout ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\valid_ctrl_inter1~0_combout ),
	.cout());
defparam \valid_ctrl_inter1~0 .lut_mask = 16'hEFFF;
defparam \valid_ctrl_inter1~0 .sum_lutc_input = "datac";

dffeas valid_ctrl_int1(
	.clk(clk),
	.d(\valid_ctrl_inter1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int1~q ),
	.prn(vcc));
defparam valid_ctrl_int1.is_wysiwyg = "true";
defparam valid_ctrl_int1.power_up = "low";

cycloneive_lcell_comb \first_data~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(\first_data~q ),
	.datac(at_source_valid_s1),
	.datad(source_ready),
	.cin(gnd),
	.combout(\first_data~0_combout ),
	.cout());
defparam \first_data~0 .lut_mask = 16'hEBBE;
defparam \first_data~0 .sum_lutc_input = "datac";

dffeas first_data(
	.clk(clk),
	.d(\first_data~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_data~q ),
	.prn(vcc));
defparam first_data.is_wysiwyg = "true";
defparam first_data.power_up = "low";

cycloneive_lcell_comb \data_select~0 (
	.dataa(at_source_valid_s1),
	.datab(\first_data~q ),
	.datac(\valid_ctrl_int1~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_select~0_combout ),
	.cout());
defparam \data_select~0 .lut_mask = 16'hFEFE;
defparam \data_select~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[7]~q ),
	.prn(vcc));
defparam \data_count_int1[7] .is_wysiwyg = "true";
defparam \data_count_int1[7] .power_up = "low";

dffeas \data_count_int[9] (
	.clk(clk),
	.d(data_count[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[9]~q ),
	.prn(vcc));
defparam \data_count_int[9] .is_wysiwyg = "true";
defparam \data_count_int[9] .power_up = "low";

dffeas \data_count_int[7] (
	.clk(clk),
	.d(data_count[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[7]~q ),
	.prn(vcc));
defparam \data_count_int[7] .is_wysiwyg = "true";
defparam \data_count_int[7] .power_up = "low";

dffeas \data_count_int[8] (
	.clk(clk),
	.d(data_count[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[8]~q ),
	.prn(vcc));
defparam \data_count_int[8] .is_wysiwyg = "true";
defparam \data_count_int[8] .power_up = "low";

dffeas \data_count_int[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[3]~q ),
	.prn(vcc));
defparam \data_count_int[3] .is_wysiwyg = "true";
defparam \data_count_int[3] .power_up = "low";

cycloneive_lcell_comb \packet_multi:count_finished~0 (
	.dataa(\data_count_int[9]~q ),
	.datab(\data_count_int[7]~q ),
	.datac(\data_count_int[8]~q ),
	.datad(\data_count_int[3]~q ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~0_combout ),
	.cout());
defparam \packet_multi:count_finished~0 .lut_mask = 16'h7FFF;
defparam \packet_multi:count_finished~0 .sum_lutc_input = "datac";

dffeas \data_count_int1[9] (
	.clk(clk),
	.d(data_count[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[9]~q ),
	.prn(vcc));
defparam \data_count_int1[9] .is_wysiwyg = "true";
defparam \data_count_int1[9] .power_up = "low";

dffeas \data_count_int1[8] (
	.clk(clk),
	.d(data_count[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[8]~q ),
	.prn(vcc));
defparam \data_count_int1[8] .is_wysiwyg = "true";
defparam \data_count_int1[8] .power_up = "low";

dffeas \data_count_int1[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[3]~q ),
	.prn(vcc));
defparam \data_count_int1[3] .is_wysiwyg = "true";
defparam \data_count_int1[3] .power_up = "low";

cycloneive_lcell_comb \packet_multi:count_finished~1 (
	.dataa(\data_count_int1[9]~q ),
	.datab(\data_count_int1[8]~q ),
	.datac(\data_count_int1[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_multi:count_finished~1_combout ),
	.cout());
defparam \packet_multi:count_finished~1 .lut_mask = 16'h7F7F;
defparam \packet_multi:count_finished~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_multi:count_finished~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int1[7]~q ),
	.datac(\packet_multi:count_finished~0_combout ),
	.datad(\packet_multi:count_finished~1_combout ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~2_combout ),
	.cout());
defparam \packet_multi:count_finished~2 .lut_mask = 16'hF7B3;
defparam \packet_multi:count_finished~2 .sum_lutc_input = "datac";

dffeas \data_count_int1[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[4]~q ),
	.prn(vcc));
defparam \data_count_int1[4] .is_wysiwyg = "true";
defparam \data_count_int1[4] .power_up = "low";

dffeas \data_count_int[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[4]~q ),
	.prn(vcc));
defparam \data_count_int[4] .is_wysiwyg = "true";
defparam \data_count_int[4] .power_up = "low";

dffeas \data_count_int[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[6]~q ),
	.prn(vcc));
defparam \data_count_int[6] .is_wysiwyg = "true";
defparam \data_count_int[6] .power_up = "low";

dffeas \data_count_int[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[5]~q ),
	.prn(vcc));
defparam \data_count_int[5] .is_wysiwyg = "true";
defparam \data_count_int[5] .power_up = "low";

dffeas \data_count_int[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[2]~q ),
	.prn(vcc));
defparam \data_count_int[2] .is_wysiwyg = "true";
defparam \data_count_int[2] .power_up = "low";

cycloneive_lcell_comb \packet_multi:count_finished~3 (
	.dataa(\data_count_int[4]~q ),
	.datab(\data_count_int[6]~q ),
	.datac(\data_count_int[5]~q ),
	.datad(\data_count_int[2]~q ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~3_combout ),
	.cout());
defparam \packet_multi:count_finished~3 .lut_mask = 16'h7FFF;
defparam \packet_multi:count_finished~3 .sum_lutc_input = "datac";

dffeas \data_count_int1[6] (
	.clk(clk),
	.d(data_count[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[6]~q ),
	.prn(vcc));
defparam \data_count_int1[6] .is_wysiwyg = "true";
defparam \data_count_int1[6] .power_up = "low";

dffeas \data_count_int1[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[5]~q ),
	.prn(vcc));
defparam \data_count_int1[5] .is_wysiwyg = "true";
defparam \data_count_int1[5] .power_up = "low";

dffeas \data_count_int1[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[2]~q ),
	.prn(vcc));
defparam \data_count_int1[2] .is_wysiwyg = "true";
defparam \data_count_int1[2] .power_up = "low";

cycloneive_lcell_comb \packet_multi:count_finished~4 (
	.dataa(\data_count_int1[6]~q ),
	.datab(\data_count_int1[5]~q ),
	.datac(\data_count_int1[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_multi:count_finished~4_combout ),
	.cout());
defparam \packet_multi:count_finished~4 .lut_mask = 16'h7F7F;
defparam \packet_multi:count_finished~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_multi:count_finished~5 (
	.dataa(\data_count_int1[4]~q ),
	.datab(\data_select~0_combout ),
	.datac(\packet_multi:count_finished~3_combout ),
	.datad(\packet_multi:count_finished~4_combout ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~5_combout ),
	.cout());
defparam \packet_multi:count_finished~5 .lut_mask = 16'hF7D5;
defparam \packet_multi:count_finished~5 .sum_lutc_input = "datac";

dffeas \data_count_int[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[0]~q ),
	.prn(vcc));
defparam \data_count_int[0] .is_wysiwyg = "true";
defparam \data_count_int[0] .power_up = "low";

dffeas \data_count_int1[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[0]~q ),
	.prn(vcc));
defparam \data_count_int1[0] .is_wysiwyg = "true";
defparam \data_count_int1[0] .power_up = "low";

dffeas \data_count_int1[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_count_int1[1]~q ),
	.prn(vcc));
defparam \data_count_int1[1] .is_wysiwyg = "true";
defparam \data_count_int1[1] .power_up = "low";

dffeas \data_count_int[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_count_int[1]~q ),
	.prn(vcc));
defparam \data_count_int[1] .is_wysiwyg = "true";
defparam \data_count_int[1] .power_up = "low";

cycloneive_lcell_comb \data_count_int_selected[1]~0 (
	.dataa(\data_count_int1[1]~q ),
	.datab(\data_count_int[1]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_count_int_selected[1]~0_combout ),
	.cout());
defparam \data_count_int_selected[1]~0 .lut_mask = 16'hAACC;
defparam \data_count_int_selected[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_multi:count_finished~6 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int[0]~q ),
	.datac(\data_count_int1[0]~q ),
	.datad(\data_count_int_selected[1]~0_combout ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~6_combout ),
	.cout());
defparam \packet_multi:count_finished~6 .lut_mask = 16'h27FF;
defparam \packet_multi:count_finished~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~0 (
	.dataa(\valid_ctrl_int~q ),
	.datab(at_source_valid_s1),
	.datac(\first_data~q ),
	.datad(\valid_ctrl_int1~q ),
	.cin(gnd),
	.combout(\at_source_valid_int~0_combout ),
	.cout());
defparam \at_source_valid_int~0 .lut_mask = 16'hFFFE;
defparam \at_source_valid_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_multi:count_finished (
	.dataa(\packet_multi:count_finished~2_combout ),
	.datab(\packet_multi:count_finished~5_combout ),
	.datac(\packet_multi:count_finished~6_combout ),
	.datad(\at_source_valid_int~0_combout ),
	.cin(gnd),
	.combout(\packet_multi:count_finished~combout ),
	.cout());
defparam \packet_multi:count_finished .lut_mask = 16'hFEFF;
defparam \packet_multi:count_finished .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\packet_multi:source_state.sop~q ),
	.datab(\packet_multi:count_finished~combout ),
	.datac(at_source_valid_s1),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(at_source_valid_s1),
	.datab(gnd),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hAAFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\packet_multi:source_state.sop~q ),
	.datab(\Selector1~0_combout ),
	.datac(source_packet_error_1),
	.datad(source_packet_error_0),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hEFFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~0 (
	.dataa(\data_count_int[3]~q ),
	.datab(\data_count_int[8]~q ),
	.datac(\data_count_int[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~0_combout ),
	.cout());
defparam \source_comb_update_2~0 .lut_mask = 16'hFEFE;
defparam \source_comb_update_2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~1 (
	.dataa(\data_count_int1[3]~q ),
	.datab(\data_count_int1[9]~q ),
	.datac(\data_count_int1[8]~q ),
	.datad(\data_count_int1[7]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~1_combout ),
	.cout());
defparam \source_comb_update_2~1 .lut_mask = 16'hFFFE;
defparam \source_comb_update_2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~2 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int[9]~q ),
	.datac(\source_comb_update_2~0_combout ),
	.datad(\source_comb_update_2~1_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~2_combout ),
	.cout());
defparam \source_comb_update_2~2 .lut_mask = 16'h27FF;
defparam \source_comb_update_2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~3 (
	.dataa(\data_count_int[6]~q ),
	.datab(\data_count_int[4]~q ),
	.datac(\data_count_int[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_comb_update_2~3_combout ),
	.cout());
defparam \source_comb_update_2~3 .lut_mask = 16'hFEFE;
defparam \source_comb_update_2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~4 (
	.dataa(\data_count_int1[6]~q ),
	.datab(\data_count_int1[5]~q ),
	.datac(\data_count_int1[4]~q ),
	.datad(\data_count_int1[2]~q ),
	.cin(gnd),
	.combout(\source_comb_update_2~4_combout ),
	.cout());
defparam \source_comb_update_2~4 .lut_mask = 16'hFFFE;
defparam \source_comb_update_2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~5 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int[5]~q ),
	.datac(\source_comb_update_2~3_combout ),
	.datad(\source_comb_update_2~4_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~5_combout ),
	.cout());
defparam \source_comb_update_2~5 .lut_mask = 16'h27FF;
defparam \source_comb_update_2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~6 (
	.dataa(\data_select~0_combout ),
	.datab(\data_count_int[0]~q ),
	.datac(\data_count_int1[0]~q ),
	.datad(\data_count_int_selected[1]~0_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~6_combout ),
	.cout());
defparam \source_comb_update_2~6 .lut_mask = 16'h27FF;
defparam \source_comb_update_2~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \source_comb_update_2~7 (
	.dataa(\at_source_valid_int~0_combout ),
	.datab(\source_comb_update_2~2_combout ),
	.datac(\source_comb_update_2~5_combout ),
	.datad(\source_comb_update_2~6_combout ),
	.cin(gnd),
	.combout(\source_comb_update_2~7_combout ),
	.cout());
defparam \source_comb_update_2~7 .lut_mask = 16'hFFFE;
defparam \source_comb_update_2~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~3 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
defparam \Selector1~3 .lut_mask = 16'hEEEE;
defparam \Selector1~3 .sum_lutc_input = "datac";

dffeas \packet_multi:source_state.st_err (
	.clk(clk),
	.d(\packet_error0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.st_err~q ),
	.prn(vcc));
defparam \packet_multi:source_state.st_err .is_wysiwyg = "true";
defparam \packet_multi:source_state.st_err .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(\packet_multi:source_state.end1~q ),
	.datad(\packet_multi:source_state.start~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFEFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(\packet_multi:source_state.st_err~q ),
	.datab(\Selector0~0_combout ),
	.datac(\source_comb_update_2~7_combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hFFF7;
defparam \Selector0~1 .sum_lutc_input = "datac";

dffeas \packet_multi:source_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.start~q ),
	.prn(vcc));
defparam \packet_multi:source_state.start .is_wysiwyg = "true";
defparam \packet_multi:source_state.start .power_up = "low";

cycloneive_lcell_comb \Selector1~4 (
	.dataa(\Selector1~3_combout ),
	.datab(\packet_multi:source_state.end1~q ),
	.datac(\packet_multi:source_state.start~q ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
defparam \Selector1~4 .lut_mask = 16'hEFFF;
defparam \Selector1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~5 (
	.dataa(\Selector1~1_combout ),
	.datab(\Selector1~2_combout ),
	.datac(\source_comb_update_2~7_combout ),
	.datad(\Selector1~4_combout ),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
defparam \Selector1~5 .lut_mask = 16'hFFFE;
defparam \Selector1~5 .sum_lutc_input = "datac";

dffeas \packet_multi:source_state.sop (
	.clk(clk),
	.d(\Selector1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.sop~q ),
	.prn(vcc));
defparam \packet_multi:source_state.sop .is_wysiwyg = "true";
defparam \packet_multi:source_state.sop .power_up = "low";

cycloneive_lcell_comb \Selector2~4 (
	.dataa(\Selector1~3_combout ),
	.datab(\packet_multi:source_state.run1~q ),
	.datac(\packet_multi:source_state.sop~q ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
defparam \Selector2~4 .lut_mask = 16'hFEFF;
defparam \Selector2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~5 (
	.dataa(\packet_multi:source_state.run1~q ),
	.datab(\packet_multi:count_finished~combout ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector2~4_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
defparam \Selector2~5 .lut_mask = 16'hFFFE;
defparam \Selector2~5 .sum_lutc_input = "datac";

dffeas \packet_multi:source_state.run1 (
	.clk(clk),
	.d(\Selector2~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.run1~q ),
	.prn(vcc));
defparam \packet_multi:source_state.run1 .is_wysiwyg = "true";
defparam \packet_multi:source_state.run1 .power_up = "low";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(\packet_multi:source_state.sop~q ),
	.datab(\packet_multi:source_state.run1~q ),
	.datac(source_packet_error_1),
	.datad(source_packet_error_0),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'hEFFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~2 (
	.dataa(\Selector3~0_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\packet_multi:count_finished~combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hEFFF;
defparam \Selector3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~1 (
	.dataa(source_packet_error_1),
	.datab(source_packet_error_0),
	.datac(source_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_source_valid_int~1_combout ),
	.cout());
defparam \at_source_valid_int~1 .lut_mask = 16'h7F7F;
defparam \at_source_valid_int~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~2 (
	.dataa(\at_source_valid_int~0_combout ),
	.datab(\packet_error0~combout ),
	.datac(at_source_valid_s1),
	.datad(\at_source_valid_int~1_combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~2_combout ),
	.cout());
defparam \at_source_valid_int~2 .lut_mask = 16'hFFFB;
defparam \at_source_valid_int~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~3 (
	.dataa(at_source_valid_s1),
	.datab(\Selector2~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\at_source_valid_int~3_combout ),
	.cout());
defparam \at_source_valid_int~3 .lut_mask = 16'hEEEE;
defparam \at_source_valid_int~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \at_source_valid_int~4 (
	.dataa(\Selector3~2_combout ),
	.datab(\Selector1~5_combout ),
	.datac(\at_source_valid_int~2_combout ),
	.datad(\at_source_valid_int~3_combout ),
	.cin(gnd),
	.combout(\at_source_valid_int~4_combout ),
	.cout());
defparam \at_source_valid_int~4 .lut_mask = 16'hFFFE;
defparam \at_source_valid_int~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\packet_error0~combout ),
	.datab(\packet_multi:source_state.end1~q ),
	.datac(\packet_multi:source_state.start~q ),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEFFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~6 (
	.dataa(at_source_valid_s1),
	.datab(source_ready),
	.datac(\packet_multi:count_finished~combout ),
	.datad(\packet_error0~combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hFBFF;
defparam \Selector2~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~1 (
	.dataa(\Selector5~0_combout ),
	.datab(\packet_multi:source_state.sop~q ),
	.datac(\packet_multi:source_state.run1~q ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

dffeas \data_int1[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[16]~q ),
	.prn(vcc));
defparam \data_int1[16] .is_wysiwyg = "true";
defparam \data_int1[16] .power_up = "low";

dffeas \data_int[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[16]~q ),
	.prn(vcc));
defparam \data_int[16] .is_wysiwyg = "true";
defparam \data_int[16] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[16]~0 (
	.dataa(\data_int1[16]~q ),
	.datab(\data_int[16]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[16]~0_combout ),
	.cout());
defparam \data_int_selected[16]~0 .lut_mask = 16'hAACC;
defparam \data_int_selected[16]~0 .sum_lutc_input = "datac";

dffeas \data_int1[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[17]~q ),
	.prn(vcc));
defparam \data_int1[17] .is_wysiwyg = "true";
defparam \data_int1[17] .power_up = "low";

dffeas \data_int[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[17]~q ),
	.prn(vcc));
defparam \data_int[17] .is_wysiwyg = "true";
defparam \data_int[17] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[17]~1 (
	.dataa(\data_int1[17]~q ),
	.datab(\data_int[17]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[17]~1_combout ),
	.cout());
defparam \data_int_selected[17]~1 .lut_mask = 16'hAACC;
defparam \data_int_selected[17]~1 .sum_lutc_input = "datac";

dffeas \data_int1[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[18]~q ),
	.prn(vcc));
defparam \data_int1[18] .is_wysiwyg = "true";
defparam \data_int1[18] .power_up = "low";

dffeas \data_int[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[18]~q ),
	.prn(vcc));
defparam \data_int[18] .is_wysiwyg = "true";
defparam \data_int[18] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[18]~2 (
	.dataa(\data_int1[18]~q ),
	.datab(\data_int[18]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[18]~2_combout ),
	.cout());
defparam \data_int_selected[18]~2 .lut_mask = 16'hAACC;
defparam \data_int_selected[18]~2 .sum_lutc_input = "datac";

dffeas \data_int1[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[19]~q ),
	.prn(vcc));
defparam \data_int1[19] .is_wysiwyg = "true";
defparam \data_int1[19] .power_up = "low";

dffeas \data_int[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[19]~q ),
	.prn(vcc));
defparam \data_int[19] .is_wysiwyg = "true";
defparam \data_int[19] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[19]~3 (
	.dataa(\data_int1[19]~q ),
	.datab(\data_int[19]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[19]~3_combout ),
	.cout());
defparam \data_int_selected[19]~3 .lut_mask = 16'hAACC;
defparam \data_int_selected[19]~3 .sum_lutc_input = "datac";

dffeas \data_int1[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[20]~q ),
	.prn(vcc));
defparam \data_int1[20] .is_wysiwyg = "true";
defparam \data_int1[20] .power_up = "low";

dffeas \data_int[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[20]~q ),
	.prn(vcc));
defparam \data_int[20] .is_wysiwyg = "true";
defparam \data_int[20] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[20]~4 (
	.dataa(\data_int1[20]~q ),
	.datab(\data_int[20]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[20]~4_combout ),
	.cout());
defparam \data_int_selected[20]~4 .lut_mask = 16'hAACC;
defparam \data_int_selected[20]~4 .sum_lutc_input = "datac";

dffeas \data_int1[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[21]~q ),
	.prn(vcc));
defparam \data_int1[21] .is_wysiwyg = "true";
defparam \data_int1[21] .power_up = "low";

dffeas \data_int[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[21]~q ),
	.prn(vcc));
defparam \data_int[21] .is_wysiwyg = "true";
defparam \data_int[21] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[21]~5 (
	.dataa(\data_int1[21]~q ),
	.datab(\data_int[21]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[21]~5_combout ),
	.cout());
defparam \data_int_selected[21]~5 .lut_mask = 16'hAACC;
defparam \data_int_selected[21]~5 .sum_lutc_input = "datac";

dffeas \data_int1[22] (
	.clk(clk),
	.d(data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[22]~q ),
	.prn(vcc));
defparam \data_int1[22] .is_wysiwyg = "true";
defparam \data_int1[22] .power_up = "low";

dffeas \data_int[22] (
	.clk(clk),
	.d(data[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[22]~q ),
	.prn(vcc));
defparam \data_int[22] .is_wysiwyg = "true";
defparam \data_int[22] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[22]~6 (
	.dataa(\data_int1[22]~q ),
	.datab(\data_int[22]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[22]~6_combout ),
	.cout());
defparam \data_int_selected[22]~6 .lut_mask = 16'hAACC;
defparam \data_int_selected[22]~6 .sum_lutc_input = "datac";

dffeas \data_int1[23] (
	.clk(clk),
	.d(data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[23]~q ),
	.prn(vcc));
defparam \data_int1[23] .is_wysiwyg = "true";
defparam \data_int1[23] .power_up = "low";

dffeas \data_int[23] (
	.clk(clk),
	.d(data[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[23]~q ),
	.prn(vcc));
defparam \data_int[23] .is_wysiwyg = "true";
defparam \data_int[23] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[23]~7 (
	.dataa(\data_int1[23]~q ),
	.datab(\data_int[23]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[23]~7_combout ),
	.cout());
defparam \data_int_selected[23]~7 .lut_mask = 16'hAACC;
defparam \data_int_selected[23]~7 .sum_lutc_input = "datac";

dffeas \data_int1[24] (
	.clk(clk),
	.d(data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[24]~q ),
	.prn(vcc));
defparam \data_int1[24] .is_wysiwyg = "true";
defparam \data_int1[24] .power_up = "low";

dffeas \data_int[24] (
	.clk(clk),
	.d(data[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[24]~q ),
	.prn(vcc));
defparam \data_int[24] .is_wysiwyg = "true";
defparam \data_int[24] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[24]~8 (
	.dataa(\data_int1[24]~q ),
	.datab(\data_int[24]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[24]~8_combout ),
	.cout());
defparam \data_int_selected[24]~8 .lut_mask = 16'hAACC;
defparam \data_int_selected[24]~8 .sum_lutc_input = "datac";

dffeas \data_int1[25] (
	.clk(clk),
	.d(data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[25]~q ),
	.prn(vcc));
defparam \data_int1[25] .is_wysiwyg = "true";
defparam \data_int1[25] .power_up = "low";

dffeas \data_int[25] (
	.clk(clk),
	.d(data[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[25]~q ),
	.prn(vcc));
defparam \data_int[25] .is_wysiwyg = "true";
defparam \data_int[25] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[25]~9 (
	.dataa(\data_int1[25]~q ),
	.datab(\data_int[25]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[25]~9_combout ),
	.cout());
defparam \data_int_selected[25]~9 .lut_mask = 16'hAACC;
defparam \data_int_selected[25]~9 .sum_lutc_input = "datac";

dffeas \data_int1[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[6]~q ),
	.prn(vcc));
defparam \data_int1[6] .is_wysiwyg = "true";
defparam \data_int1[6] .power_up = "low";

dffeas \data_int[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[6]~q ),
	.prn(vcc));
defparam \data_int[6] .is_wysiwyg = "true";
defparam \data_int[6] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[6]~10 (
	.dataa(\data_int1[6]~q ),
	.datab(\data_int[6]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[6]~10_combout ),
	.cout());
defparam \data_int_selected[6]~10 .lut_mask = 16'hAACC;
defparam \data_int_selected[6]~10 .sum_lutc_input = "datac";

dffeas \data_int1[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[7]~q ),
	.prn(vcc));
defparam \data_int1[7] .is_wysiwyg = "true";
defparam \data_int1[7] .power_up = "low";

dffeas \data_int[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[7]~q ),
	.prn(vcc));
defparam \data_int[7] .is_wysiwyg = "true";
defparam \data_int[7] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[7]~11 (
	.dataa(\data_int1[7]~q ),
	.datab(\data_int[7]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[7]~11_combout ),
	.cout());
defparam \data_int_selected[7]~11 .lut_mask = 16'hAACC;
defparam \data_int_selected[7]~11 .sum_lutc_input = "datac";

dffeas \data_int1[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[8]~q ),
	.prn(vcc));
defparam \data_int1[8] .is_wysiwyg = "true";
defparam \data_int1[8] .power_up = "low";

dffeas \data_int[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[8]~q ),
	.prn(vcc));
defparam \data_int[8] .is_wysiwyg = "true";
defparam \data_int[8] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[8]~12 (
	.dataa(\data_int1[8]~q ),
	.datab(\data_int[8]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[8]~12_combout ),
	.cout());
defparam \data_int_selected[8]~12 .lut_mask = 16'hAACC;
defparam \data_int_selected[8]~12 .sum_lutc_input = "datac";

dffeas \data_int1[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[9]~q ),
	.prn(vcc));
defparam \data_int1[9] .is_wysiwyg = "true";
defparam \data_int1[9] .power_up = "low";

dffeas \data_int[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[9]~q ),
	.prn(vcc));
defparam \data_int[9] .is_wysiwyg = "true";
defparam \data_int[9] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[9]~13 (
	.dataa(\data_int1[9]~q ),
	.datab(\data_int[9]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[9]~13_combout ),
	.cout());
defparam \data_int_selected[9]~13 .lut_mask = 16'hAACC;
defparam \data_int_selected[9]~13 .sum_lutc_input = "datac";

dffeas \data_int1[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[10]~q ),
	.prn(vcc));
defparam \data_int1[10] .is_wysiwyg = "true";
defparam \data_int1[10] .power_up = "low";

dffeas \data_int[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[10]~q ),
	.prn(vcc));
defparam \data_int[10] .is_wysiwyg = "true";
defparam \data_int[10] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[10]~14 (
	.dataa(\data_int1[10]~q ),
	.datab(\data_int[10]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[10]~14_combout ),
	.cout());
defparam \data_int_selected[10]~14 .lut_mask = 16'hAACC;
defparam \data_int_selected[10]~14 .sum_lutc_input = "datac";

dffeas \data_int1[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[11]~q ),
	.prn(vcc));
defparam \data_int1[11] .is_wysiwyg = "true";
defparam \data_int1[11] .power_up = "low";

dffeas \data_int[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[11]~q ),
	.prn(vcc));
defparam \data_int[11] .is_wysiwyg = "true";
defparam \data_int[11] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[11]~15 (
	.dataa(\data_int1[11]~q ),
	.datab(\data_int[11]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[11]~15_combout ),
	.cout());
defparam \data_int_selected[11]~15 .lut_mask = 16'hAACC;
defparam \data_int_selected[11]~15 .sum_lutc_input = "datac";

dffeas \data_int1[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[12]~q ),
	.prn(vcc));
defparam \data_int1[12] .is_wysiwyg = "true";
defparam \data_int1[12] .power_up = "low";

dffeas \data_int[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[12]~q ),
	.prn(vcc));
defparam \data_int[12] .is_wysiwyg = "true";
defparam \data_int[12] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[12]~16 (
	.dataa(\data_int1[12]~q ),
	.datab(\data_int[12]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[12]~16_combout ),
	.cout());
defparam \data_int_selected[12]~16 .lut_mask = 16'hAACC;
defparam \data_int_selected[12]~16 .sum_lutc_input = "datac";

dffeas \data_int1[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[13]~q ),
	.prn(vcc));
defparam \data_int1[13] .is_wysiwyg = "true";
defparam \data_int1[13] .power_up = "low";

dffeas \data_int[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[13]~q ),
	.prn(vcc));
defparam \data_int[13] .is_wysiwyg = "true";
defparam \data_int[13] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[13]~17 (
	.dataa(\data_int1[13]~q ),
	.datab(\data_int[13]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[13]~17_combout ),
	.cout());
defparam \data_int_selected[13]~17 .lut_mask = 16'hAACC;
defparam \data_int_selected[13]~17 .sum_lutc_input = "datac";

dffeas \data_int1[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[14]~q ),
	.prn(vcc));
defparam \data_int1[14] .is_wysiwyg = "true";
defparam \data_int1[14] .power_up = "low";

dffeas \data_int[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[14]~q ),
	.prn(vcc));
defparam \data_int[14] .is_wysiwyg = "true";
defparam \data_int[14] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[14]~18 (
	.dataa(\data_int1[14]~q ),
	.datab(\data_int[14]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[14]~18_combout ),
	.cout());
defparam \data_int_selected[14]~18 .lut_mask = 16'hAACC;
defparam \data_int_selected[14]~18 .sum_lutc_input = "datac";

dffeas \data_int1[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[15]~q ),
	.prn(vcc));
defparam \data_int1[15] .is_wysiwyg = "true";
defparam \data_int1[15] .power_up = "low";

dffeas \data_int[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[15]~q ),
	.prn(vcc));
defparam \data_int[15] .is_wysiwyg = "true";
defparam \data_int[15] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[15]~19 (
	.dataa(\data_int1[15]~q ),
	.datab(\data_int[15]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[15]~19_combout ),
	.cout());
defparam \data_int_selected[15]~19 .lut_mask = 16'hAACC;
defparam \data_int_selected[15]~19 .sum_lutc_input = "datac";

dffeas \data_int1[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[0]~q ),
	.prn(vcc));
defparam \data_int1[0] .is_wysiwyg = "true";
defparam \data_int1[0] .power_up = "low";

dffeas \data_int[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[0]~q ),
	.prn(vcc));
defparam \data_int[0] .is_wysiwyg = "true";
defparam \data_int[0] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[0]~20 (
	.dataa(\data_int1[0]~q ),
	.datab(\data_int[0]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[0]~20_combout ),
	.cout());
defparam \data_int_selected[0]~20 .lut_mask = 16'hAACC;
defparam \data_int_selected[0]~20 .sum_lutc_input = "datac";

dffeas \data_int1[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[1]~q ),
	.prn(vcc));
defparam \data_int1[1] .is_wysiwyg = "true";
defparam \data_int1[1] .power_up = "low";

dffeas \data_int[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[1]~q ),
	.prn(vcc));
defparam \data_int[1] .is_wysiwyg = "true";
defparam \data_int[1] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[1]~21 (
	.dataa(\data_int1[1]~q ),
	.datab(\data_int[1]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[1]~21_combout ),
	.cout());
defparam \data_int_selected[1]~21 .lut_mask = 16'hAACC;
defparam \data_int_selected[1]~21 .sum_lutc_input = "datac";

dffeas \data_int1[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[2]~q ),
	.prn(vcc));
defparam \data_int1[2] .is_wysiwyg = "true";
defparam \data_int1[2] .power_up = "low";

dffeas \data_int[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[2]~q ),
	.prn(vcc));
defparam \data_int[2] .is_wysiwyg = "true";
defparam \data_int[2] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[2]~22 (
	.dataa(\data_int1[2]~q ),
	.datab(\data_int[2]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[2]~22_combout ),
	.cout());
defparam \data_int_selected[2]~22 .lut_mask = 16'hAACC;
defparam \data_int_selected[2]~22 .sum_lutc_input = "datac";

dffeas \data_int1[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[3]~q ),
	.prn(vcc));
defparam \data_int1[3] .is_wysiwyg = "true";
defparam \data_int1[3] .power_up = "low";

dffeas \data_int[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[3]~q ),
	.prn(vcc));
defparam \data_int[3] .is_wysiwyg = "true";
defparam \data_int[3] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[3]~23 (
	.dataa(\data_int1[3]~q ),
	.datab(\data_int[3]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[3]~23_combout ),
	.cout());
defparam \data_int_selected[3]~23 .lut_mask = 16'hAACC;
defparam \data_int_selected[3]~23 .sum_lutc_input = "datac";

dffeas \data_int1[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[4]~q ),
	.prn(vcc));
defparam \data_int1[4] .is_wysiwyg = "true";
defparam \data_int1[4] .power_up = "low";

dffeas \data_int[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[4]~q ),
	.prn(vcc));
defparam \data_int[4] .is_wysiwyg = "true";
defparam \data_int[4] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[4]~24 (
	.dataa(\data_int1[4]~q ),
	.datab(\data_int[4]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[4]~24_combout ),
	.cout());
defparam \data_int_selected[4]~24 .lut_mask = 16'hAACC;
defparam \data_int_selected[4]~24 .sum_lutc_input = "datac";

dffeas \data_int1[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~0_combout ),
	.q(\data_int1[5]~q ),
	.prn(vcc));
defparam \data_int1[5] .is_wysiwyg = "true";
defparam \data_int1[5] .power_up = "low";

dffeas \data_int[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~1_combout ),
	.q(\data_int[5]~q ),
	.prn(vcc));
defparam \data_int[5] .is_wysiwyg = "true";
defparam \data_int[5] .power_up = "low";

cycloneive_lcell_comb \data_int_selected[5]~25 (
	.dataa(\data_int1[5]~q ),
	.datab(\data_int[5]~q ),
	.datac(gnd),
	.datad(\data_select~0_combout ),
	.cin(gnd),
	.combout(\data_int_selected[5]~25_combout ),
	.cout());
defparam \data_int_selected[5]~25 .lut_mask = 16'hAACC;
defparam \data_int_selected[5]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\valid_ctrl_int1~q ),
	.datab(\first_data~q ),
	.datac(source_ready),
	.datad(at_source_valid_s1),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFBF;
defparam \Mux0~0 .sum_lutc_input = "datac";

endmodule
