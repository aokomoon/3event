module DDS
#(

)
(
    input       wire        sys_clk     ,
    input       wire        sys_rst     ,
    
    
);





































endmodule 

